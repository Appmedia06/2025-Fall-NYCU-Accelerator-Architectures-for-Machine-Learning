// Copyright 2021 The CFU-Playground Authors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.



module Cfu (
  input               cmd_valid,
  output reg          cmd_ready,
  input      [9:0]    cmd_payload_function_id,
  input      [31:0]   cmd_payload_inputs_0,
  input      [31:0]   cmd_payload_inputs_1,
  output reg          rsp_valid,
  input               rsp_ready,
  output reg [31:0]   rsp_payload_outputs_0,
  input               reset,
  input               clk
);

wire data_en = cmd_valid && cmd_ready;

reg [31:0] input_data0;
always @(posedge clk) begin
  if ( reset ) begin
    input_data0 <= 32'd0;
  end
  else if ( data_en ) begin
    input_data0 <= cmd_payload_inputs_0;
  end
end


wire [9:0]  recip_addr = input_data0[30:21];
reg  [31:0] recip_out;
always @( * ) begin
    case ( recip_addr )
      10'h000: recip_out = 32'h7FFFFFFF; // x = 0.0000, f(x) = 1.0000
      10'h001: recip_out = 32'h7FE007FE; // x = 0.0010, f(x) = 0.9990
      10'h002: recip_out = 32'h7FC01FF0; // x = 0.0020, f(x) = 0.9981
      10'h003: recip_out = 32'h7FA047CA; // x = 0.0029, f(x) = 0.9971
      10'h004: recip_out = 32'h7F807F80; // x = 0.0039, f(x) = 0.9961
      10'h005: recip_out = 32'h7F60C707; // x = 0.0049, f(x) = 0.9951
      10'h006: recip_out = 32'h7F411E53; // x = 0.0059, f(x) = 0.9942
      10'h007: recip_out = 32'h7F218557; // x = 0.0068, f(x) = 0.9932
      10'h008: recip_out = 32'h7F01FC08; // x = 0.0078, f(x) = 0.9922
      10'h009: recip_out = 32'h7EE2825B; // x = 0.0088, f(x) = 0.9913
      10'h00A: recip_out = 32'h7EC31843; // x = 0.0098, f(x) = 0.9903
      10'h00B: recip_out = 32'h7EA3BDB6; // x = 0.0107, f(x) = 0.9894
      10'h00C: recip_out = 32'h7E8472A8; // x = 0.0117, f(x) = 0.9884
      10'h00D: recip_out = 32'h7E65370D; // x = 0.0127, f(x) = 0.9875
      10'h00E: recip_out = 32'h7E460ADA; // x = 0.0137, f(x) = 0.9865
      10'h00F: recip_out = 32'h7E26EE03; // x = 0.0146, f(x) = 0.9856
      10'h010: recip_out = 32'h7E07E07E; // x = 0.0156, f(x) = 0.9846
      10'h011: recip_out = 32'h7DE8E23E; // x = 0.0166, f(x) = 0.9837
      10'h012: recip_out = 32'h7DC9F339; // x = 0.0176, f(x) = 0.9827
      10'h013: recip_out = 32'h7DAB1364; // x = 0.0186, f(x) = 0.9818
      10'h014: recip_out = 32'h7D8C42B3; // x = 0.0195, f(x) = 0.9808
      10'h015: recip_out = 32'h7D6D811A; // x = 0.0205, f(x) = 0.9799
      10'h016: recip_out = 32'h7D4ECE90; // x = 0.0215, f(x) = 0.9790
      10'h017: recip_out = 32'h7D302B09; // x = 0.0225, f(x) = 0.9780
      10'h018: recip_out = 32'h7D119679; // x = 0.0234, f(x) = 0.9771
      10'h019: recip_out = 32'h7CF310D7; // x = 0.0244, f(x) = 0.9762
      10'h01A: recip_out = 32'h7CD49A16; // x = 0.0254, f(x) = 0.9752
      10'h01B: recip_out = 32'h7CB6322D; // x = 0.0264, f(x) = 0.9743
      10'h01C: recip_out = 32'h7C97D911; // x = 0.0273, f(x) = 0.9734
      10'h01D: recip_out = 32'h7C798EB5; // x = 0.0283, f(x) = 0.9725
      10'h01E: recip_out = 32'h7C5B5311; // x = 0.0293, f(x) = 0.9715
      10'h01F: recip_out = 32'h7C3D2619; // x = 0.0303, f(x) = 0.9706
      10'h020: recip_out = 32'h7C1F07C2; // x = 0.0312, f(x) = 0.9697
      10'h021: recip_out = 32'h7C00F802; // x = 0.0322, f(x) = 0.9688
      10'h022: recip_out = 32'h7BE2F6CE; // x = 0.0332, f(x) = 0.9679
      10'h023: recip_out = 32'h7BC5041C; // x = 0.0342, f(x) = 0.9669
      10'h024: recip_out = 32'h7BA71FE1; // x = 0.0352, f(x) = 0.9660
      10'h025: recip_out = 32'h7B894A13; // x = 0.0361, f(x) = 0.9651
      10'h026: recip_out = 32'h7B6B82A7; // x = 0.0371, f(x) = 0.9642
      10'h027: recip_out = 32'h7B4DC993; // x = 0.0381, f(x) = 0.9633
      10'h028: recip_out = 32'h7B301ECC; // x = 0.0391, f(x) = 0.9624
      10'h029: recip_out = 32'h7B128249; // x = 0.0400, f(x) = 0.9615
      10'h02A: recip_out = 32'h7AF4F3FE; // x = 0.0410, f(x) = 0.9606
      10'h02B: recip_out = 32'h7AD773E2; // x = 0.0420, f(x) = 0.9597
      10'h02C: recip_out = 32'h7ABA01EB; // x = 0.0430, f(x) = 0.9588
      10'h02D: recip_out = 32'h7A9C9E0E; // x = 0.0439, f(x) = 0.9579
      10'h02E: recip_out = 32'h7A7F4841; // x = 0.0449, f(x) = 0.9570
      10'h02F: recip_out = 32'h7A62007A; // x = 0.0459, f(x) = 0.9561
      10'h030: recip_out = 32'h7A44C6B0; // x = 0.0469, f(x) = 0.9552
      10'h031: recip_out = 32'h7A279AD7; // x = 0.0479, f(x) = 0.9543
      10'h032: recip_out = 32'h7A0A7CE7; // x = 0.0488, f(x) = 0.9534
      10'h033: recip_out = 32'h79ED6CD4; // x = 0.0498, f(x) = 0.9526
      10'h034: recip_out = 32'h79D06A96; // x = 0.0508, f(x) = 0.9517
      10'h035: recip_out = 32'h79B37623; // x = 0.0518, f(x) = 0.9508
      10'h036: recip_out = 32'h79968F70; // x = 0.0527, f(x) = 0.9499
      10'h037: recip_out = 32'h7979B673; // x = 0.0537, f(x) = 0.9490
      10'h038: recip_out = 32'h795CEB24; // x = 0.0547, f(x) = 0.9481
      10'h039: recip_out = 32'h79402D78; // x = 0.0557, f(x) = 0.9473
      10'h03A: recip_out = 32'h79237D66; // x = 0.0566, f(x) = 0.9464
      10'h03B: recip_out = 32'h7906DAE3; // x = 0.0576, f(x) = 0.9455
      10'h03C: recip_out = 32'h78EA45E7; // x = 0.0586, f(x) = 0.9446
      10'h03D: recip_out = 32'h78CDBE68; // x = 0.0596, f(x) = 0.9438
      10'h03E: recip_out = 32'h78B1445C; // x = 0.0605, f(x) = 0.9429
      10'h03F: recip_out = 32'h7894D7BA; // x = 0.0615, f(x) = 0.9420
      10'h040: recip_out = 32'h78787878; // x = 0.0625, f(x) = 0.9412
      10'h041: recip_out = 32'h785C268E; // x = 0.0635, f(x) = 0.9403
      10'h042: recip_out = 32'h783FE1F0; // x = 0.0645, f(x) = 0.9394
      10'h043: recip_out = 32'h7823AA97; // x = 0.0654, f(x) = 0.9386
      10'h044: recip_out = 32'h78078078; // x = 0.0664, f(x) = 0.9377
      10'h045: recip_out = 32'h77EB638B; // x = 0.0674, f(x) = 0.9369
      10'h046: recip_out = 32'h77CF53C6; // x = 0.0684, f(x) = 0.9360
      10'h047: recip_out = 32'h77B35120; // x = 0.0693, f(x) = 0.9352
      10'h048: recip_out = 32'h77975B90; // x = 0.0703, f(x) = 0.9343
      10'h049: recip_out = 32'h777B730C; // x = 0.0713, f(x) = 0.9335
      10'h04A: recip_out = 32'h775F978C; // x = 0.0723, f(x) = 0.9326
      10'h04B: recip_out = 32'h7743C907; // x = 0.0732, f(x) = 0.9318
      10'h04C: recip_out = 32'h77280773; // x = 0.0742, f(x) = 0.9309
      10'h04D: recip_out = 32'h770C52C7; // x = 0.0752, f(x) = 0.9301
      10'h04E: recip_out = 32'h76F0AAFA; // x = 0.0762, f(x) = 0.9292
      10'h04F: recip_out = 32'h76D51004; // x = 0.0771, f(x) = 0.9284
      10'h050: recip_out = 32'h76B981DB; // x = 0.0781, f(x) = 0.9275
      10'h051: recip_out = 32'h769E0077; // x = 0.0791, f(x) = 0.9267
      10'h052: recip_out = 32'h76828BCE; // x = 0.0801, f(x) = 0.9259
      10'h053: recip_out = 32'h766723D8; // x = 0.0811, f(x) = 0.9250
      10'h054: recip_out = 32'h764BC88C; // x = 0.0820, f(x) = 0.9242
      10'h055: recip_out = 32'h763079E2; // x = 0.0830, f(x) = 0.9234
      10'h056: recip_out = 32'h761537D0; // x = 0.0840, f(x) = 0.9225
      10'h057: recip_out = 32'h75FA024E; // x = 0.0850, f(x) = 0.9217
      10'h058: recip_out = 32'h75DED953; // x = 0.0859, f(x) = 0.9209
      10'h059: recip_out = 32'h75C3BCD6; // x = 0.0869, f(x) = 0.9200
      10'h05A: recip_out = 32'h75A8ACD0; // x = 0.0879, f(x) = 0.9192
      10'h05B: recip_out = 32'h758DA936; // x = 0.0889, f(x) = 0.9184
      10'h05C: recip_out = 32'h7572B202; // x = 0.0898, f(x) = 0.9176
      10'h05D: recip_out = 32'h7557C729; // x = 0.0908, f(x) = 0.9167
      10'h05E: recip_out = 32'h753CE8A5; // x = 0.0918, f(x) = 0.9159
      10'h05F: recip_out = 32'h7522166C; // x = 0.0928, f(x) = 0.9151
      10'h060: recip_out = 32'h75075075; // x = 0.0938, f(x) = 0.9143
      10'h061: recip_out = 32'h74EC96B9; // x = 0.0947, f(x) = 0.9135
      10'h062: recip_out = 32'h74D1E92F; // x = 0.0957, f(x) = 0.9127
      10'h063: recip_out = 32'h74B747CF; // x = 0.0967, f(x) = 0.9118
      10'h064: recip_out = 32'h749CB290; // x = 0.0977, f(x) = 0.9110
      10'h065: recip_out = 32'h7482296A; // x = 0.0986, f(x) = 0.9102
      10'h066: recip_out = 32'h7467AC55; // x = 0.0996, f(x) = 0.9094
      10'h067: recip_out = 32'h744D3B49; // x = 0.1006, f(x) = 0.9086
      10'h068: recip_out = 32'h7432D63E; // x = 0.1016, f(x) = 0.9078
      10'h069: recip_out = 32'h74187D2A; // x = 0.1025, f(x) = 0.9070
      10'h06A: recip_out = 32'h73FE3007; // x = 0.1035, f(x) = 0.9062
      10'h06B: recip_out = 32'h73E3EECC; // x = 0.1045, f(x) = 0.9054
      10'h06C: recip_out = 32'h73C9B971; // x = 0.1055, f(x) = 0.9046
      10'h06D: recip_out = 32'h73AF8FEE; // x = 0.1064, f(x) = 0.9038
      10'h06E: recip_out = 32'h7395723B; // x = 0.1074, f(x) = 0.9030
      10'h06F: recip_out = 32'h737B604F; // x = 0.1084, f(x) = 0.9022
      10'h070: recip_out = 32'h73615A24; // x = 0.1094, f(x) = 0.9014
      10'h071: recip_out = 32'h73475FB1; // x = 0.1104, f(x) = 0.9006
      10'h072: recip_out = 32'h732D70EE; // x = 0.1113, f(x) = 0.8998
      10'h073: recip_out = 32'h73138DD3; // x = 0.1123, f(x) = 0.8990
      10'h074: recip_out = 32'h72F9B658; // x = 0.1133, f(x) = 0.8982
      10'h075: recip_out = 32'h72DFEA76; // x = 0.1143, f(x) = 0.8975
      10'h076: recip_out = 32'h72C62A25; // x = 0.1152, f(x) = 0.8967
      10'h077: recip_out = 32'h72AC755D; // x = 0.1162, f(x) = 0.8959
      10'h078: recip_out = 32'h7292CC15; // x = 0.1172, f(x) = 0.8951
      10'h079: recip_out = 32'h72792E48; // x = 0.1182, f(x) = 0.8943
      10'h07A: recip_out = 32'h725F9BEC; // x = 0.1191, f(x) = 0.8935
      10'h07B: recip_out = 32'h724614FB; // x = 0.1201, f(x) = 0.8928
      10'h07C: recip_out = 32'h722C996C; // x = 0.1211, f(x) = 0.8920
      10'h07D: recip_out = 32'h72132938; // x = 0.1221, f(x) = 0.8912
      10'h07E: recip_out = 32'h71F9C457; // x = 0.1230, f(x) = 0.8904
      10'h07F: recip_out = 32'h71E06AC2; // x = 0.1240, f(x) = 0.8897
      10'h080: recip_out = 32'h71C71C72; // x = 0.1250, f(x) = 0.8889
      10'h081: recip_out = 32'h71ADD95E; // x = 0.1260, f(x) = 0.8881
      10'h082: recip_out = 32'h7194A17F; // x = 0.1270, f(x) = 0.8873
      10'h083: recip_out = 32'h717B74CF; // x = 0.1279, f(x) = 0.8866
      10'h084: recip_out = 32'h71625344; // x = 0.1289, f(x) = 0.8858
      10'h085: recip_out = 32'h71493CD9; // x = 0.1299, f(x) = 0.8850
      10'h086: recip_out = 32'h71303185; // x = 0.1309, f(x) = 0.8843
      10'h087: recip_out = 32'h71173142; // x = 0.1318, f(x) = 0.8835
      10'h088: recip_out = 32'h70FE3C07; // x = 0.1328, f(x) = 0.8828
      10'h089: recip_out = 32'h70E551CE; // x = 0.1338, f(x) = 0.8820
      10'h08A: recip_out = 32'h70CC7290; // x = 0.1348, f(x) = 0.8812
      10'h08B: recip_out = 32'h70B39E44; // x = 0.1357, f(x) = 0.8805
      10'h08C: recip_out = 32'h709AD4E5; // x = 0.1367, f(x) = 0.8797
      10'h08D: recip_out = 32'h7082166A; // x = 0.1377, f(x) = 0.8790
      10'h08E: recip_out = 32'h706962CD; // x = 0.1387, f(x) = 0.8782
      10'h08F: recip_out = 32'h7050BA06; // x = 0.1396, f(x) = 0.8775
      10'h090: recip_out = 32'h70381C0E; // x = 0.1406, f(x) = 0.8767
      10'h091: recip_out = 32'h701F88DE; // x = 0.1416, f(x) = 0.8760
      10'h092: recip_out = 32'h70070070; // x = 0.1426, f(x) = 0.8752
      10'h093: recip_out = 32'h6FEE82BC; // x = 0.1436, f(x) = 0.8745
      10'h094: recip_out = 32'h6FD60FBA; // x = 0.1445, f(x) = 0.8737
      10'h095: recip_out = 32'h6FBDA765; // x = 0.1455, f(x) = 0.8730
      10'h096: recip_out = 32'h6FA549B4; // x = 0.1465, f(x) = 0.8722
      10'h097: recip_out = 32'h6F8CF6A2; // x = 0.1475, f(x) = 0.8715
      10'h098: recip_out = 32'h6F74AE26; // x = 0.1484, f(x) = 0.8707
      10'h099: recip_out = 32'h6F5C703B; // x = 0.1494, f(x) = 0.8700
      10'h09A: recip_out = 32'h6F443CD9; // x = 0.1504, f(x) = 0.8693
      10'h09B: recip_out = 32'h6F2C13FA; // x = 0.1514, f(x) = 0.8685
      10'h09C: recip_out = 32'h6F13F596; // x = 0.1523, f(x) = 0.8678
      10'h09D: recip_out = 32'h6EFBE1A7; // x = 0.1533, f(x) = 0.8671
      10'h09E: recip_out = 32'h6EE3D826; // x = 0.1543, f(x) = 0.8663
      10'h09F: recip_out = 32'h6ECBD90C; // x = 0.1553, f(x) = 0.8656
      10'h0A0: recip_out = 32'h6EB3E453; // x = 0.1562, f(x) = 0.8649
      10'h0A1: recip_out = 32'h6E9BF9F3; // x = 0.1572, f(x) = 0.8641
      10'h0A2: recip_out = 32'h6E8419E7; // x = 0.1582, f(x) = 0.8634
      10'h0A3: recip_out = 32'h6E6C4427; // x = 0.1592, f(x) = 0.8627
      10'h0A4: recip_out = 32'h6E5478AC; // x = 0.1602, f(x) = 0.8620
      10'h0A5: recip_out = 32'h6E3CB771; // x = 0.1611, f(x) = 0.8612
      10'h0A6: recip_out = 32'h6E25006E; // x = 0.1621, f(x) = 0.8605
      10'h0A7: recip_out = 32'h6E0D539D; // x = 0.1631, f(x) = 0.8598
      10'h0A8: recip_out = 32'h6DF5B0F7; // x = 0.1641, f(x) = 0.8591
      10'h0A9: recip_out = 32'h6DDE1876; // x = 0.1650, f(x) = 0.8583
      10'h0AA: recip_out = 32'h6DC68A14; // x = 0.1660, f(x) = 0.8576
      10'h0AB: recip_out = 32'h6DAF05C9; // x = 0.1670, f(x) = 0.8569
      10'h0AC: recip_out = 32'h6D978B8F; // x = 0.1680, f(x) = 0.8562
      10'h0AD: recip_out = 32'h6D801B60; // x = 0.1689, f(x) = 0.8555
      10'h0AE: recip_out = 32'h6D68B535; // x = 0.1699, f(x) = 0.8548
      10'h0AF: recip_out = 32'h6D515909; // x = 0.1709, f(x) = 0.8540
      10'h0B0: recip_out = 32'h6D3A06D4; // x = 0.1719, f(x) = 0.8533
      10'h0B1: recip_out = 32'h6D22BE90; // x = 0.1729, f(x) = 0.8526
      10'h0B2: recip_out = 32'h6D0B8037; // x = 0.1738, f(x) = 0.8519
      10'h0B3: recip_out = 32'h6CF44BC2; // x = 0.1748, f(x) = 0.8512
      10'h0B4: recip_out = 32'h6CDD212B; // x = 0.1758, f(x) = 0.8505
      10'h0B5: recip_out = 32'h6CC6006D; // x = 0.1768, f(x) = 0.8498
      10'h0B6: recip_out = 32'h6CAEE980; // x = 0.1777, f(x) = 0.8491
      10'h0B7: recip_out = 32'h6C97DC5E; // x = 0.1787, f(x) = 0.8484
      10'h0B8: recip_out = 32'h6C80D902; // x = 0.1797, f(x) = 0.8477
      10'h0B9: recip_out = 32'h6C69DF64; // x = 0.1807, f(x) = 0.8470
      10'h0BA: recip_out = 32'h6C52EF7F; // x = 0.1816, f(x) = 0.8463
      10'h0BB: recip_out = 32'h6C3C094D; // x = 0.1826, f(x) = 0.8456
      10'h0BC: recip_out = 32'h6C252CC7; // x = 0.1836, f(x) = 0.8449
      10'h0BD: recip_out = 32'h6C0E59E8; // x = 0.1846, f(x) = 0.8442
      10'h0BE: recip_out = 32'h6BF790A9; // x = 0.1855, f(x) = 0.8435
      10'h0BF: recip_out = 32'h6BE0D104; // x = 0.1865, f(x) = 0.8428
      10'h0C0: recip_out = 32'h6BCA1AF3; // x = 0.1875, f(x) = 0.8421
      10'h0C1: recip_out = 32'h6BB36E6F; // x = 0.1885, f(x) = 0.8414
      10'h0C2: recip_out = 32'h6B9CCB74; // x = 0.1895, f(x) = 0.8407
      10'h0C3: recip_out = 32'h6B8631FB; // x = 0.1904, f(x) = 0.8400
      10'h0C4: recip_out = 32'h6B6FA1FE; // x = 0.1914, f(x) = 0.8393
      10'h0C5: recip_out = 32'h6B591B77; // x = 0.1924, f(x) = 0.8387
      10'h0C6: recip_out = 32'h6B429E60; // x = 0.1934, f(x) = 0.8380
      10'h0C7: recip_out = 32'h6B2C2AB4; // x = 0.1943, f(x) = 0.8373
      10'h0C8: recip_out = 32'h6B15C06B; // x = 0.1953, f(x) = 0.8366
      10'h0C9: recip_out = 32'h6AFF5F81; // x = 0.1963, f(x) = 0.8359
      10'h0CA: recip_out = 32'h6AE907EF; // x = 0.1973, f(x) = 0.8352
      10'h0CB: recip_out = 32'h6AD2B9B0; // x = 0.1982, f(x) = 0.8346
      10'h0CC: recip_out = 32'h6ABC74BE; // x = 0.1992, f(x) = 0.8339
      10'h0CD: recip_out = 32'h6AA63913; // x = 0.2002, f(x) = 0.8332
      10'h0CE: recip_out = 32'h6A9006A9; // x = 0.2012, f(x) = 0.8325
      10'h0CF: recip_out = 32'h6A79DD7A; // x = 0.2021, f(x) = 0.8318
      10'h0D0: recip_out = 32'h6A63BD82; // x = 0.2031, f(x) = 0.8312
      10'h0D1: recip_out = 32'h6A4DA6B9; // x = 0.2041, f(x) = 0.8305
      10'h0D2: recip_out = 32'h6A37991A; // x = 0.2051, f(x) = 0.8298
      10'h0D3: recip_out = 32'h6A2194A0; // x = 0.2061, f(x) = 0.8291
      10'h0D4: recip_out = 32'h6A0B9945; // x = 0.2070, f(x) = 0.8285
      10'h0D5: recip_out = 32'h69F5A703; // x = 0.2080, f(x) = 0.8278
      10'h0D6: recip_out = 32'h69DFBDD4; // x = 0.2090, f(x) = 0.8271
      10'h0D7: recip_out = 32'h69C9DDB4; // x = 0.2100, f(x) = 0.8265
      10'h0D8: recip_out = 32'h69B4069B; // x = 0.2109, f(x) = 0.8258
      10'h0D9: recip_out = 32'h699E3886; // x = 0.2119, f(x) = 0.8251
      10'h0DA: recip_out = 32'h6988736D; // x = 0.2129, f(x) = 0.8245
      10'h0DB: recip_out = 32'h6972B74C; // x = 0.2139, f(x) = 0.8238
      10'h0DC: recip_out = 32'h695D041E; // x = 0.2148, f(x) = 0.8232
      10'h0DD: recip_out = 32'h694759DB; // x = 0.2158, f(x) = 0.8225
      10'h0DE: recip_out = 32'h6931B880; // x = 0.2168, f(x) = 0.8218
      10'h0DF: recip_out = 32'h691C2007; // x = 0.2178, f(x) = 0.8212
      10'h0E0: recip_out = 32'h69069069; // x = 0.2188, f(x) = 0.8205
      10'h0E1: recip_out = 32'h68F109A2; // x = 0.2197, f(x) = 0.8199
      10'h0E2: recip_out = 32'h68DB8BAC; // x = 0.2207, f(x) = 0.8192
      10'h0E3: recip_out = 32'h68C61683; // x = 0.2217, f(x) = 0.8185
      10'h0E4: recip_out = 32'h68B0AA1F; // x = 0.2227, f(x) = 0.8179
      10'h0E5: recip_out = 32'h689B467D; // x = 0.2236, f(x) = 0.8172
      10'h0E6: recip_out = 32'h6885EB96; // x = 0.2246, f(x) = 0.8166
      10'h0E7: recip_out = 32'h68709965; // x = 0.2256, f(x) = 0.8159
      10'h0E8: recip_out = 32'h685B4FE6; // x = 0.2266, f(x) = 0.8153
      10'h0E9: recip_out = 32'h68460F12; // x = 0.2275, f(x) = 0.8146
      10'h0EA: recip_out = 32'h6830D6E5; // x = 0.2285, f(x) = 0.8140
      10'h0EB: recip_out = 32'h681BA758; // x = 0.2295, f(x) = 0.8133
      10'h0EC: recip_out = 32'h68068068; // x = 0.2305, f(x) = 0.8127
      10'h0ED: recip_out = 32'h67F1620E; // x = 0.2314, f(x) = 0.8121
      10'h0EE: recip_out = 32'h67DC4C46; // x = 0.2324, f(x) = 0.8114
      10'h0EF: recip_out = 32'h67C73F0A; // x = 0.2334, f(x) = 0.8108
      10'h0F0: recip_out = 32'h67B23A54; // x = 0.2344, f(x) = 0.8101
      10'h0F1: recip_out = 32'h679D3E21; // x = 0.2354, f(x) = 0.8095
      10'h0F2: recip_out = 32'h67884A6A; // x = 0.2363, f(x) = 0.8088
      10'h0F3: recip_out = 32'h67735F2B; // x = 0.2373, f(x) = 0.8082
      10'h0F4: recip_out = 32'h675E7C5E; // x = 0.2383, f(x) = 0.8076
      10'h0F5: recip_out = 32'h6749A1FE; // x = 0.2393, f(x) = 0.8069
      10'h0F6: recip_out = 32'h6734D006; // x = 0.2402, f(x) = 0.8063
      10'h0F7: recip_out = 32'h67200672; // x = 0.2412, f(x) = 0.8057
      10'h0F8: recip_out = 32'h670B453C; // x = 0.2422, f(x) = 0.8050
      10'h0F9: recip_out = 32'h66F68C5E; // x = 0.2432, f(x) = 0.8044
      10'h0FA: recip_out = 32'h66E1DBD5; // x = 0.2441, f(x) = 0.8038
      10'h0FB: recip_out = 32'h66CD339A; // x = 0.2451, f(x) = 0.8031
      10'h0FC: recip_out = 32'h66B893A9; // x = 0.2461, f(x) = 0.8025
      10'h0FD: recip_out = 32'h66A3FBFE; // x = 0.2471, f(x) = 0.8019
      10'h0FE: recip_out = 32'h668F6C92; // x = 0.2480, f(x) = 0.8013
      10'h0FF: recip_out = 32'h667AE561; // x = 0.2490, f(x) = 0.8006
      10'h100: recip_out = 32'h66666666; // x = 0.2500, f(x) = 0.8000
      10'h101: recip_out = 32'h6651EF9D; // x = 0.2510, f(x) = 0.7994
      10'h102: recip_out = 32'h663D8100; // x = 0.2520, f(x) = 0.7988
      10'h103: recip_out = 32'h66291A8A; // x = 0.2529, f(x) = 0.7981
      10'h104: recip_out = 32'h6614BC36; // x = 0.2539, f(x) = 0.7975
      10'h105: recip_out = 32'h66006600; // x = 0.2549, f(x) = 0.7969
      10'h106: recip_out = 32'h65EC17E3; // x = 0.2559, f(x) = 0.7963
      10'h107: recip_out = 32'h65D7D1DA; // x = 0.2568, f(x) = 0.7956
      10'h108: recip_out = 32'h65C393E0; // x = 0.2578, f(x) = 0.7950
      10'h109: recip_out = 32'h65AF5DF1; // x = 0.2588, f(x) = 0.7944
      10'h10A: recip_out = 32'h659B3006; // x = 0.2598, f(x) = 0.7938
      10'h10B: recip_out = 32'h65870A1D; // x = 0.2607, f(x) = 0.7932
      10'h10C: recip_out = 32'h6572EC30; // x = 0.2617, f(x) = 0.7926
      10'h10D: recip_out = 32'h655ED639; // x = 0.2627, f(x) = 0.7920
      10'h10E: recip_out = 32'h654AC836; // x = 0.2637, f(x) = 0.7913
      10'h10F: recip_out = 32'h6536C220; // x = 0.2646, f(x) = 0.7907
      10'h110: recip_out = 32'h6522C3F3; // x = 0.2656, f(x) = 0.7901
      10'h111: recip_out = 32'h650ECDAB; // x = 0.2666, f(x) = 0.7895
      10'h112: recip_out = 32'h64FADF43; // x = 0.2676, f(x) = 0.7889
      10'h113: recip_out = 32'h64E6F8B5; // x = 0.2686, f(x) = 0.7883
      10'h114: recip_out = 32'h64D319FE; // x = 0.2695, f(x) = 0.7877
      10'h115: recip_out = 32'h64BF4319; // x = 0.2705, f(x) = 0.7871
      10'h116: recip_out = 32'h64AB7402; // x = 0.2715, f(x) = 0.7865
      10'h117: recip_out = 32'h6497ACB2; // x = 0.2725, f(x) = 0.7859
      10'h118: recip_out = 32'h6483ED27; // x = 0.2734, f(x) = 0.7853
      10'h119: recip_out = 32'h6470355C; // x = 0.2744, f(x) = 0.7847
      10'h11A: recip_out = 32'h645C854B; // x = 0.2754, f(x) = 0.7841
      10'h11B: recip_out = 32'h6448DCF1; // x = 0.2764, f(x) = 0.7835
      10'h11C: recip_out = 32'h64353C48; // x = 0.2773, f(x) = 0.7829
      10'h11D: recip_out = 32'h6421A34D; // x = 0.2783, f(x) = 0.7823
      10'h11E: recip_out = 32'h640E11FB; // x = 0.2793, f(x) = 0.7817
      10'h11F: recip_out = 32'h63FA884D; // x = 0.2803, f(x) = 0.7811
      10'h120: recip_out = 32'h63E7063E; // x = 0.2812, f(x) = 0.7805
      10'h121: recip_out = 32'h63D38BCC; // x = 0.2822, f(x) = 0.7799
      10'h122: recip_out = 32'h63C018F0; // x = 0.2832, f(x) = 0.7793
      10'h123: recip_out = 32'h63ACADA7; // x = 0.2842, f(x) = 0.7787
      10'h124: recip_out = 32'h639949EC; // x = 0.2852, f(x) = 0.7781
      10'h125: recip_out = 32'h6385EDBA; // x = 0.2861, f(x) = 0.7775
      10'h126: recip_out = 32'h6372990E; // x = 0.2871, f(x) = 0.7769
      10'h127: recip_out = 32'h635F4BE3; // x = 0.2881, f(x) = 0.7763
      10'h128: recip_out = 32'h634C0635; // x = 0.2891, f(x) = 0.7758
      10'h129: recip_out = 32'h6338C7FE; // x = 0.2900, f(x) = 0.7752
      10'h12A: recip_out = 32'h6325913C; // x = 0.2910, f(x) = 0.7746
      10'h12B: recip_out = 32'h631261E9; // x = 0.2920, f(x) = 0.7740
      10'h12C: recip_out = 32'h62FF3A02; // x = 0.2930, f(x) = 0.7734
      10'h12D: recip_out = 32'h62EC1981; // x = 0.2939, f(x) = 0.7728
      10'h12E: recip_out = 32'h62D90063; // x = 0.2949, f(x) = 0.7722
      10'h12F: recip_out = 32'h62C5EEA3; // x = 0.2959, f(x) = 0.7717
      10'h130: recip_out = 32'h62B2E43E; // x = 0.2969, f(x) = 0.7711
      10'h131: recip_out = 32'h629FE12E; // x = 0.2979, f(x) = 0.7705
      10'h132: recip_out = 32'h628CE570; // x = 0.2988, f(x) = 0.7699
      10'h133: recip_out = 32'h6279F0FF; // x = 0.2998, f(x) = 0.7693
      10'h134: recip_out = 32'h626703D8; // x = 0.3008, f(x) = 0.7688
      10'h135: recip_out = 32'h62541DF6; // x = 0.3018, f(x) = 0.7682
      10'h136: recip_out = 32'h62413F54; // x = 0.3027, f(x) = 0.7676
      10'h137: recip_out = 32'h622E67EF; // x = 0.3037, f(x) = 0.7670
      10'h138: recip_out = 32'h621B97C3; // x = 0.3047, f(x) = 0.7665
      10'h139: recip_out = 32'h6208CECB; // x = 0.3057, f(x) = 0.7659
      10'h13A: recip_out = 32'h61F60D03; // x = 0.3066, f(x) = 0.7653
      10'h13B: recip_out = 32'h61E35267; // x = 0.3076, f(x) = 0.7647
      10'h13C: recip_out = 32'h61D09EF3; // x = 0.3086, f(x) = 0.7642
      10'h13D: recip_out = 32'h61BDF2A3; // x = 0.3096, f(x) = 0.7636
      10'h13E: recip_out = 32'h61AB4D73; // x = 0.3105, f(x) = 0.7630
      10'h13F: recip_out = 32'h6198AF5E; // x = 0.3115, f(x) = 0.7625
      10'h140: recip_out = 32'h61861862; // x = 0.3125, f(x) = 0.7619
      10'h141: recip_out = 32'h61738878; // x = 0.3135, f(x) = 0.7613
      10'h142: recip_out = 32'h6160FF9F; // x = 0.3145, f(x) = 0.7608
      10'h143: recip_out = 32'h614E7DD0; // x = 0.3154, f(x) = 0.7602
      10'h144: recip_out = 32'h613C030A; // x = 0.3164, f(x) = 0.7596
      10'h145: recip_out = 32'h61298F47; // x = 0.3174, f(x) = 0.7591
      10'h146: recip_out = 32'h61172283; // x = 0.3184, f(x) = 0.7585
      10'h147: recip_out = 32'h6104BCBB; // x = 0.3193, f(x) = 0.7580
      10'h148: recip_out = 32'h60F25DEB; // x = 0.3203, f(x) = 0.7574
      10'h149: recip_out = 32'h60E0060E; // x = 0.3213, f(x) = 0.7568
      10'h14A: recip_out = 32'h60CDB521; // x = 0.3223, f(x) = 0.7563
      10'h14B: recip_out = 32'h60BB6B20; // x = 0.3232, f(x) = 0.7557
      10'h14C: recip_out = 32'h60A92806; // x = 0.3242, f(x) = 0.7552
      10'h14D: recip_out = 32'h6096EBD0; // x = 0.3252, f(x) = 0.7546
      10'h14E: recip_out = 32'h6084B67B; // x = 0.3262, f(x) = 0.7541
      10'h14F: recip_out = 32'h60728802; // x = 0.3271, f(x) = 0.7535
      10'h150: recip_out = 32'h60606060; // x = 0.3281, f(x) = 0.7529
      10'h151: recip_out = 32'h604E3F94; // x = 0.3291, f(x) = 0.7524
      10'h152: recip_out = 32'h603C2597; // x = 0.3301, f(x) = 0.7518
      10'h153: recip_out = 32'h602A1268; // x = 0.3311, f(x) = 0.7513
      10'h154: recip_out = 32'h60180602; // x = 0.3320, f(x) = 0.7507
      10'h155: recip_out = 32'h60060060; // x = 0.3330, f(x) = 0.7502
      10'h156: recip_out = 32'h5FF40180; // x = 0.3340, f(x) = 0.7496
      10'h157: recip_out = 32'h5FE2095D; // x = 0.3350, f(x) = 0.7491
      10'h158: recip_out = 32'h5FD017F4; // x = 0.3359, f(x) = 0.7485
      10'h159: recip_out = 32'h5FBE2D41; // x = 0.3369, f(x) = 0.7480
      10'h15A: recip_out = 32'h5FAC4940; // x = 0.3379, f(x) = 0.7474
      10'h15B: recip_out = 32'h5F9A6BED; // x = 0.3389, f(x) = 0.7469
      10'h15C: recip_out = 32'h5F889545; // x = 0.3398, f(x) = 0.7464
      10'h15D: recip_out = 32'h5F76C544; // x = 0.3408, f(x) = 0.7458
      10'h15E: recip_out = 32'h5F64FBE7; // x = 0.3418, f(x) = 0.7453
      10'h15F: recip_out = 32'h5F533928; // x = 0.3428, f(x) = 0.7447
      10'h160: recip_out = 32'h5F417D06; // x = 0.3438, f(x) = 0.7442
      10'h161: recip_out = 32'h5F2FC77C; // x = 0.3447, f(x) = 0.7436
      10'h162: recip_out = 32'h5F1E1886; // x = 0.3457, f(x) = 0.7431
      10'h163: recip_out = 32'h5F0C7021; // x = 0.3467, f(x) = 0.7426
      10'h164: recip_out = 32'h5EFACE49; // x = 0.3477, f(x) = 0.7420
      10'h165: recip_out = 32'h5EE932FA; // x = 0.3486, f(x) = 0.7415
      10'h166: recip_out = 32'h5ED79E32; // x = 0.3496, f(x) = 0.7410
      10'h167: recip_out = 32'h5EC60FEB; // x = 0.3506, f(x) = 0.7404
      10'h168: recip_out = 32'h5EB48824; // x = 0.3516, f(x) = 0.7399
      10'h169: recip_out = 32'h5EA306D7; // x = 0.3525, f(x) = 0.7394
      10'h16A: recip_out = 32'h5E918C01; // x = 0.3535, f(x) = 0.7388
      10'h16B: recip_out = 32'h5E8017A0; // x = 0.3545, f(x) = 0.7383
      10'h16C: recip_out = 32'h5E6EA9AF; // x = 0.3555, f(x) = 0.7378
      10'h16D: recip_out = 32'h5E5D422A; // x = 0.3564, f(x) = 0.7372
      10'h16E: recip_out = 32'h5E4BE10F; // x = 0.3574, f(x) = 0.7367
      10'h16F: recip_out = 32'h5E3A8659; // x = 0.3584, f(x) = 0.7362
      10'h170: recip_out = 32'h5E293206; // x = 0.3594, f(x) = 0.7356
      10'h171: recip_out = 32'h5E17E411; // x = 0.3604, f(x) = 0.7351
      10'h172: recip_out = 32'h5E069C77; // x = 0.3613, f(x) = 0.7346
      10'h173: recip_out = 32'h5DF55B35; // x = 0.3623, f(x) = 0.7341
      10'h174: recip_out = 32'h5DE42046; // x = 0.3633, f(x) = 0.7335
      10'h175: recip_out = 32'h5DD2EBA9; // x = 0.3643, f(x) = 0.7330
      10'h176: recip_out = 32'h5DC1BD58; // x = 0.3652, f(x) = 0.7325
      10'h177: recip_out = 32'h5DB09551; // x = 0.3662, f(x) = 0.7320
      10'h178: recip_out = 32'h5D9F7391; // x = 0.3672, f(x) = 0.7314
      10'h179: recip_out = 32'h5D8E5813; // x = 0.3682, f(x) = 0.7309
      10'h17A: recip_out = 32'h5D7D42D5; // x = 0.3691, f(x) = 0.7304
      10'h17B: recip_out = 32'h5D6C33D2; // x = 0.3701, f(x) = 0.7299
      10'h17C: recip_out = 32'h5D5B2B08; // x = 0.3711, f(x) = 0.7293
      10'h17D: recip_out = 32'h5D4A2873; // x = 0.3721, f(x) = 0.7288
      10'h17E: recip_out = 32'h5D392C10; // x = 0.3730, f(x) = 0.7283
      10'h17F: recip_out = 32'h5D2835DB; // x = 0.3740, f(x) = 0.7278
      10'h180: recip_out = 32'h5D1745D1; // x = 0.3750, f(x) = 0.7273
      10'h181: recip_out = 32'h5D065BEF; // x = 0.3760, f(x) = 0.7268
      10'h182: recip_out = 32'h5CF57831; // x = 0.3770, f(x) = 0.7262
      10'h183: recip_out = 32'h5CE49A94; // x = 0.3779, f(x) = 0.7257
      10'h184: recip_out = 32'h5CD3C315; // x = 0.3789, f(x) = 0.7252
      10'h185: recip_out = 32'h5CC2F1B0; // x = 0.3799, f(x) = 0.7247
      10'h186: recip_out = 32'h5CB22662; // x = 0.3809, f(x) = 0.7242
      10'h187: recip_out = 32'h5CA16127; // x = 0.3818, f(x) = 0.7237
      10'h188: recip_out = 32'h5C90A1FD; // x = 0.3828, f(x) = 0.7232
      10'h189: recip_out = 32'h5C7FE8E0; // x = 0.3838, f(x) = 0.7227
      10'h18A: recip_out = 32'h5C6F35CD; // x = 0.3848, f(x) = 0.7221
      10'h18B: recip_out = 32'h5C5E88C0; // x = 0.3857, f(x) = 0.7216
      10'h18C: recip_out = 32'h5C4DE1B6; // x = 0.3867, f(x) = 0.7211
      10'h18D: recip_out = 32'h5C3D40AD; // x = 0.3877, f(x) = 0.7206
      10'h18E: recip_out = 32'h5C2CA5A0; // x = 0.3887, f(x) = 0.7201
      10'h18F: recip_out = 32'h5C1C108D; // x = 0.3896, f(x) = 0.7196
      10'h190: recip_out = 32'h5C0B8170; // x = 0.3906, f(x) = 0.7191
      10'h191: recip_out = 32'h5BFAF846; // x = 0.3916, f(x) = 0.7186
      10'h192: recip_out = 32'h5BEA750D; // x = 0.3926, f(x) = 0.7181
      10'h193: recip_out = 32'h5BD9F7BF; // x = 0.3936, f(x) = 0.7176
      10'h194: recip_out = 32'h5BC9805C; // x = 0.3945, f(x) = 0.7171
      10'h195: recip_out = 32'h5BB90EDE; // x = 0.3955, f(x) = 0.7166
      10'h196: recip_out = 32'h5BA8A344; // x = 0.3965, f(x) = 0.7161
      10'h197: recip_out = 32'h5B983D8A; // x = 0.3975, f(x) = 0.7156
      10'h198: recip_out = 32'h5B87DDAD; // x = 0.3984, f(x) = 0.7151
      10'h199: recip_out = 32'h5B7783AA; // x = 0.3994, f(x) = 0.7146
      10'h19A: recip_out = 32'h5B672F7D; // x = 0.4004, f(x) = 0.7141
      10'h19B: recip_out = 32'h5B56E123; // x = 0.4014, f(x) = 0.7136
      10'h19C: recip_out = 32'h5B46989A; // x = 0.4023, f(x) = 0.7131
      10'h19D: recip_out = 32'h5B3655DE; // x = 0.4033, f(x) = 0.7126
      10'h19E: recip_out = 32'h5B2618EC; // x = 0.4043, f(x) = 0.7121
      10'h19F: recip_out = 32'h5B15E1C2; // x = 0.4053, f(x) = 0.7116
      10'h1A0: recip_out = 32'h5B05B05B; // x = 0.4062, f(x) = 0.7111
      10'h1A1: recip_out = 32'h5AF584B5; // x = 0.4072, f(x) = 0.7106
      10'h1A2: recip_out = 32'h5AE55ECD; // x = 0.4082, f(x) = 0.7101
      10'h1A3: recip_out = 32'h5AD53EA0; // x = 0.4092, f(x) = 0.7096
      10'h1A4: recip_out = 32'h5AC5242B; // x = 0.4102, f(x) = 0.7091
      10'h1A5: recip_out = 32'h5AB50F6A; // x = 0.4111, f(x) = 0.7087
      10'h1A6: recip_out = 32'h5AA5005B; // x = 0.4121, f(x) = 0.7082
      10'h1A7: recip_out = 32'h5A94F6FA; // x = 0.4131, f(x) = 0.7077
      10'h1A8: recip_out = 32'h5A84F345; // x = 0.4141, f(x) = 0.7072
      10'h1A9: recip_out = 32'h5A74F539; // x = 0.4150, f(x) = 0.7067
      10'h1AA: recip_out = 32'h5A64FCD2; // x = 0.4160, f(x) = 0.7062
      10'h1AB: recip_out = 32'h5A550A0E; // x = 0.4170, f(x) = 0.7057
      10'h1AC: recip_out = 32'h5A451CEA; // x = 0.4180, f(x) = 0.7052
      10'h1AD: recip_out = 32'h5A353562; // x = 0.4189, f(x) = 0.7047
      10'h1AE: recip_out = 32'h5A255375; // x = 0.4199, f(x) = 0.7043
      10'h1AF: recip_out = 32'h5A15771D; // x = 0.4209, f(x) = 0.7038
      10'h1B0: recip_out = 32'h5A05A05A; // x = 0.4219, f(x) = 0.7033
      10'h1B1: recip_out = 32'h59F5CF28; // x = 0.4229, f(x) = 0.7028
      10'h1B2: recip_out = 32'h59E60383; // x = 0.4238, f(x) = 0.7023
      10'h1B3: recip_out = 32'h59D63D69; // x = 0.4248, f(x) = 0.7019
      10'h1B4: recip_out = 32'h59C67CD8; // x = 0.4258, f(x) = 0.7014
      10'h1B5: recip_out = 32'h59B6C1CC; // x = 0.4268, f(x) = 0.7009
      10'h1B6: recip_out = 32'h59A70C42; // x = 0.4277, f(x) = 0.7004
      10'h1B7: recip_out = 32'h59975C37; // x = 0.4287, f(x) = 0.6999
      10'h1B8: recip_out = 32'h5987B1A9; // x = 0.4297, f(x) = 0.6995
      10'h1B9: recip_out = 32'h59780C95; // x = 0.4307, f(x) = 0.6990
      10'h1BA: recip_out = 32'h59686CF7; // x = 0.4316, f(x) = 0.6985
      10'h1BB: recip_out = 32'h5958D2CE; // x = 0.4326, f(x) = 0.6980
      10'h1BC: recip_out = 32'h59493E15; // x = 0.4336, f(x) = 0.6975
      10'h1BD: recip_out = 32'h5939AECA; // x = 0.4346, f(x) = 0.6971
      10'h1BE: recip_out = 32'h592A24EB; // x = 0.4355, f(x) = 0.6966
      10'h1BF: recip_out = 32'h591AA075; // x = 0.4365, f(x) = 0.6961
      10'h1C0: recip_out = 32'h590B2164; // x = 0.4375, f(x) = 0.6957
      10'h1C1: recip_out = 32'h58FBA7B6; // x = 0.4385, f(x) = 0.6952
      10'h1C2: recip_out = 32'h58EC3369; // x = 0.4395, f(x) = 0.6947
      10'h1C3: recip_out = 32'h58DCC478; // x = 0.4404, f(x) = 0.6942
      10'h1C4: recip_out = 32'h58CD5AE2; // x = 0.4414, f(x) = 0.6938
      10'h1C5: recip_out = 32'h58BDF6A4; // x = 0.4424, f(x) = 0.6933
      10'h1C6: recip_out = 32'h58AE97BB; // x = 0.4434, f(x) = 0.6928
      10'h1C7: recip_out = 32'h589F3E24; // x = 0.4443, f(x) = 0.6924
      10'h1C8: recip_out = 32'h588FE9DC; // x = 0.4453, f(x) = 0.6919
      10'h1C9: recip_out = 32'h58809AE1; // x = 0.4463, f(x) = 0.6914
      10'h1CA: recip_out = 32'h58715130; // x = 0.4473, f(x) = 0.6910
      10'h1CB: recip_out = 32'h58620CC6; // x = 0.4482, f(x) = 0.6905
      10'h1CC: recip_out = 32'h5852CDA1; // x = 0.4492, f(x) = 0.6900
      10'h1CD: recip_out = 32'h584393BD; // x = 0.4502, f(x) = 0.6896
      10'h1CE: recip_out = 32'h58345F18; // x = 0.4512, f(x) = 0.6891
      10'h1CF: recip_out = 32'h58252FB0; // x = 0.4521, f(x) = 0.6886
      10'h1D0: recip_out = 32'h58160581; // x = 0.4531, f(x) = 0.6882
      10'h1D1: recip_out = 32'h5806E08A; // x = 0.4541, f(x) = 0.6877
      10'h1D2: recip_out = 32'h57F7C0C6; // x = 0.4551, f(x) = 0.6872
      10'h1D3: recip_out = 32'h57E8A634; // x = 0.4561, f(x) = 0.6868
      10'h1D4: recip_out = 32'h57D990D1; // x = 0.4570, f(x) = 0.6863
      10'h1D5: recip_out = 32'h57CA809A; // x = 0.4580, f(x) = 0.6859
      10'h1D6: recip_out = 32'h57BB758C; // x = 0.4590, f(x) = 0.6854
      10'h1D7: recip_out = 32'h57AC6FA6; // x = 0.4600, f(x) = 0.6849
      10'h1D8: recip_out = 32'h579D6EE3; // x = 0.4609, f(x) = 0.6845
      10'h1D9: recip_out = 32'h578E7343; // x = 0.4619, f(x) = 0.6840
      10'h1DA: recip_out = 32'h577F7CC1; // x = 0.4629, f(x) = 0.6836
      10'h1DB: recip_out = 32'h57708B5B; // x = 0.4639, f(x) = 0.6831
      10'h1DC: recip_out = 32'h57619F10; // x = 0.4648, f(x) = 0.6827
      10'h1DD: recip_out = 32'h5752B7DB; // x = 0.4658, f(x) = 0.6822
      10'h1DE: recip_out = 32'h5743D5BB; // x = 0.4668, f(x) = 0.6818
      10'h1DF: recip_out = 32'h5734F8AD; // x = 0.4678, f(x) = 0.6813
      10'h1E0: recip_out = 32'h572620AE; // x = 0.4688, f(x) = 0.6809
      10'h1E1: recip_out = 32'h57174DBC; // x = 0.4697, f(x) = 0.6804
      10'h1E2: recip_out = 32'h57087FD4; // x = 0.4707, f(x) = 0.6799
      10'h1E3: recip_out = 32'h56F9B6F4; // x = 0.4717, f(x) = 0.6795
      10'h1E4: recip_out = 32'h56EAF319; // x = 0.4727, f(x) = 0.6790
      10'h1E5: recip_out = 32'h56DC3440; // x = 0.4736, f(x) = 0.6786
      10'h1E6: recip_out = 32'h56CD7A68; // x = 0.4746, f(x) = 0.6781
      10'h1E7: recip_out = 32'h56BEC58C; // x = 0.4756, f(x) = 0.6777
      10'h1E8: recip_out = 32'h56B015AC; // x = 0.4766, f(x) = 0.6772
      10'h1E9: recip_out = 32'h56A16AC4; // x = 0.4775, f(x) = 0.6768
      10'h1EA: recip_out = 32'h5692C4D2; // x = 0.4785, f(x) = 0.6764
      10'h1EB: recip_out = 32'h568423D3; // x = 0.4795, f(x) = 0.6759
      10'h1EC: recip_out = 32'h567587C5; // x = 0.4805, f(x) = 0.6755
      10'h1ED: recip_out = 32'h5666F0A5; // x = 0.4814, f(x) = 0.6750
      10'h1EE: recip_out = 32'h56585E71; // x = 0.4824, f(x) = 0.6746
      10'h1EF: recip_out = 32'h5649D126; // x = 0.4834, f(x) = 0.6741
      10'h1F0: recip_out = 32'h563B48C2; // x = 0.4844, f(x) = 0.6737
      10'h1F1: recip_out = 32'h562CC542; // x = 0.4854, f(x) = 0.6732
      10'h1F2: recip_out = 32'h561E46A5; // x = 0.4863, f(x) = 0.6728
      10'h1F3: recip_out = 32'h560FCCE7; // x = 0.4873, f(x) = 0.6724
      10'h1F4: recip_out = 32'h56015805; // x = 0.4883, f(x) = 0.6719
      10'h1F5: recip_out = 32'h55F2E7FF; // x = 0.4893, f(x) = 0.6715
      10'h1F6: recip_out = 32'h55E47CD0; // x = 0.4902, f(x) = 0.6710
      10'h1F7: recip_out = 32'h55D61677; // x = 0.4912, f(x) = 0.6706
      10'h1F8: recip_out = 32'h55C7B4F1; // x = 0.4922, f(x) = 0.6702
      10'h1F9: recip_out = 32'h55B9583C; // x = 0.4932, f(x) = 0.6697
      10'h1FA: recip_out = 32'h55AB0056; // x = 0.4941, f(x) = 0.6693
      10'h1FB: recip_out = 32'h559CAD3B; // x = 0.4951, f(x) = 0.6688
      10'h1FC: recip_out = 32'h558E5EEA; // x = 0.4961, f(x) = 0.6684
      10'h1FD: recip_out = 32'h55801560; // x = 0.4971, f(x) = 0.6680
      10'h1FE: recip_out = 32'h5571D09B; // x = 0.4980, f(x) = 0.6675
      10'h1FF: recip_out = 32'h55639098; // x = 0.4990, f(x) = 0.6671
      10'h200: recip_out = 32'h55555555; // x = 0.5000, f(x) = 0.6667
      10'h201: recip_out = 32'h55471ED0; // x = 0.5010, f(x) = 0.6662
      10'h202: recip_out = 32'h5538ED06; // x = 0.5020, f(x) = 0.6658
      10'h203: recip_out = 32'h552ABFF5; // x = 0.5029, f(x) = 0.6654
      10'h204: recip_out = 32'h551C979B; // x = 0.5039, f(x) = 0.6649
      10'h205: recip_out = 32'h550E73F5; // x = 0.5049, f(x) = 0.6645
      10'h206: recip_out = 32'h55005500; // x = 0.5059, f(x) = 0.6641
      10'h207: recip_out = 32'h54F23ABB; // x = 0.5068, f(x) = 0.6636
      10'h208: recip_out = 32'h54E42524; // x = 0.5078, f(x) = 0.6632
      10'h209: recip_out = 32'h54D61437; // x = 0.5088, f(x) = 0.6628
      10'h20A: recip_out = 32'h54C807F3; // x = 0.5098, f(x) = 0.6624
      10'h20B: recip_out = 32'h54BA0055; // x = 0.5107, f(x) = 0.6619
      10'h20C: recip_out = 32'h54ABFD5B; // x = 0.5117, f(x) = 0.6615
      10'h20D: recip_out = 32'h549DFF02; // x = 0.5127, f(x) = 0.6611
      10'h20E: recip_out = 32'h54900549; // x = 0.5137, f(x) = 0.6606
      10'h20F: recip_out = 32'h5482102D; // x = 0.5146, f(x) = 0.6602
      10'h210: recip_out = 32'h54741FAC; // x = 0.5156, f(x) = 0.6598
      10'h211: recip_out = 32'h546633C3; // x = 0.5166, f(x) = 0.6594
      10'h212: recip_out = 32'h54584C70; // x = 0.5176, f(x) = 0.6589
      10'h213: recip_out = 32'h544A69B1; // x = 0.5186, f(x) = 0.6585
      10'h214: recip_out = 32'h543C8B84; // x = 0.5195, f(x) = 0.6581
      10'h215: recip_out = 32'h542EB1E7; // x = 0.5205, f(x) = 0.6577
      10'h216: recip_out = 32'h5420DCD6; // x = 0.5215, f(x) = 0.6573
      10'h217: recip_out = 32'h54130C51; // x = 0.5225, f(x) = 0.6568
      10'h218: recip_out = 32'h54054054; // x = 0.5234, f(x) = 0.6564
      10'h219: recip_out = 32'h53F778DE; // x = 0.5244, f(x) = 0.6560
      10'h21A: recip_out = 32'h53E9B5EC; // x = 0.5254, f(x) = 0.6556
      10'h21B: recip_out = 32'h53DBF77C; // x = 0.5264, f(x) = 0.6552
      10'h21C: recip_out = 32'h53CE3D8B; // x = 0.5273, f(x) = 0.6547
      10'h21D: recip_out = 32'h53C08819; // x = 0.5283, f(x) = 0.6543
      10'h21E: recip_out = 32'h53B2D722; // x = 0.5293, f(x) = 0.6539
      10'h21F: recip_out = 32'h53A52AA4; // x = 0.5303, f(x) = 0.6535
      10'h220: recip_out = 32'h5397829D; // x = 0.5312, f(x) = 0.6531
      10'h221: recip_out = 32'h5389DF0B; // x = 0.5322, f(x) = 0.6526
      10'h222: recip_out = 32'h537C3FEB; // x = 0.5332, f(x) = 0.6522
      10'h223: recip_out = 32'h536EA53C; // x = 0.5342, f(x) = 0.6518
      10'h224: recip_out = 32'h53610EFB; // x = 0.5352, f(x) = 0.6514
      10'h225: recip_out = 32'h53537D27; // x = 0.5361, f(x) = 0.6510
      10'h226: recip_out = 32'h5345EFBC; // x = 0.5371, f(x) = 0.6506
      10'h227: recip_out = 32'h533866BA; // x = 0.5381, f(x) = 0.6502
      10'h228: recip_out = 32'h532AE21D; // x = 0.5391, f(x) = 0.6497
      10'h229: recip_out = 32'h531D61E3; // x = 0.5400, f(x) = 0.6493
      10'h22A: recip_out = 32'h530FE60B; // x = 0.5410, f(x) = 0.6489
      10'h22B: recip_out = 32'h53026E92; // x = 0.5420, f(x) = 0.6485
      10'h22C: recip_out = 32'h52F4FB77; // x = 0.5430, f(x) = 0.6481
      10'h22D: recip_out = 32'h52E78CB6; // x = 0.5439, f(x) = 0.6477
      10'h22E: recip_out = 32'h52DA224E; // x = 0.5449, f(x) = 0.6473
      10'h22F: recip_out = 32'h52CCBC3D; // x = 0.5459, f(x) = 0.6469
      10'h230: recip_out = 32'h52BF5A81; // x = 0.5469, f(x) = 0.6465
      10'h231: recip_out = 32'h52B1FD18; // x = 0.5479, f(x) = 0.6461
      10'h232: recip_out = 32'h52A4A3FF; // x = 0.5488, f(x) = 0.6456
      10'h233: recip_out = 32'h52974F34; // x = 0.5498, f(x) = 0.6452
      10'h234: recip_out = 32'h5289FEB6; // x = 0.5508, f(x) = 0.6448
      10'h235: recip_out = 32'h527CB282; // x = 0.5518, f(x) = 0.6444
      10'h236: recip_out = 32'h526F6A96; // x = 0.5527, f(x) = 0.6440
      10'h237: recip_out = 32'h526226F0; // x = 0.5537, f(x) = 0.6436
      10'h238: recip_out = 32'h5254E78F; // x = 0.5547, f(x) = 0.6432
      10'h239: recip_out = 32'h5247AC6F; // x = 0.5557, f(x) = 0.6428
      10'h23A: recip_out = 32'h523A7590; // x = 0.5566, f(x) = 0.6424
      10'h23B: recip_out = 32'h522D42EE; // x = 0.5576, f(x) = 0.6420
      10'h23C: recip_out = 32'h52201488; // x = 0.5586, f(x) = 0.6416
      10'h23D: recip_out = 32'h5212EA5C; // x = 0.5596, f(x) = 0.6412
      10'h23E: recip_out = 32'h5205C468; // x = 0.5605, f(x) = 0.6408
      10'h23F: recip_out = 32'h51F8A2A9; // x = 0.5615, f(x) = 0.6404
      10'h240: recip_out = 32'h51EB851F; // x = 0.5625, f(x) = 0.6400
      10'h241: recip_out = 32'h51DE6BC6; // x = 0.5635, f(x) = 0.6396
      10'h242: recip_out = 32'h51D1569D; // x = 0.5645, f(x) = 0.6392
      10'h243: recip_out = 32'h51C445A1; // x = 0.5654, f(x) = 0.6388
      10'h244: recip_out = 32'h51B738D1; // x = 0.5664, f(x) = 0.6384
      10'h245: recip_out = 32'h51AA302B; // x = 0.5674, f(x) = 0.6380
      10'h246: recip_out = 32'h519D2BAD; // x = 0.5684, f(x) = 0.6376
      10'h247: recip_out = 32'h51902B55; // x = 0.5693, f(x) = 0.6372
      10'h248: recip_out = 32'h51832F20; // x = 0.5703, f(x) = 0.6368
      10'h249: recip_out = 32'h5176370D; // x = 0.5713, f(x) = 0.6364
      10'h24A: recip_out = 32'h5169431A; // x = 0.5723, f(x) = 0.6360
      10'h24B: recip_out = 32'h515C5344; // x = 0.5732, f(x) = 0.6356
      10'h24C: recip_out = 32'h514F678B; // x = 0.5742, f(x) = 0.6352
      10'h24D: recip_out = 32'h51427FEC; // x = 0.5752, f(x) = 0.6348
      10'h24E: recip_out = 32'h51359C64; // x = 0.5762, f(x) = 0.6344
      10'h24F: recip_out = 32'h5128BCF3; // x = 0.5771, f(x) = 0.6341
      10'h250: recip_out = 32'h511BE196; // x = 0.5781, f(x) = 0.6337
      10'h251: recip_out = 32'h510F0A4A; // x = 0.5791, f(x) = 0.6333
      10'h252: recip_out = 32'h51023710; // x = 0.5801, f(x) = 0.6329
      10'h253: recip_out = 32'h50F567E3; // x = 0.5811, f(x) = 0.6325
      10'h254: recip_out = 32'h50E89CC3; // x = 0.5820, f(x) = 0.6321
      10'h255: recip_out = 32'h50DBD5AD; // x = 0.5830, f(x) = 0.6317
      10'h256: recip_out = 32'h50CF12A0; // x = 0.5840, f(x) = 0.6313
      10'h257: recip_out = 32'h50C25399; // x = 0.5850, f(x) = 0.6309
      10'h258: recip_out = 32'h50B59897; // x = 0.5859, f(x) = 0.6305
      10'h259: recip_out = 32'h50A8E198; // x = 0.5869, f(x) = 0.6302
      10'h25A: recip_out = 32'h509C2E9A; // x = 0.5879, f(x) = 0.6298
      10'h25B: recip_out = 32'h508F7F9B; // x = 0.5889, f(x) = 0.6294
      10'h25C: recip_out = 32'h5082D499; // x = 0.5898, f(x) = 0.6290
      10'h25D: recip_out = 32'h50762D93; // x = 0.5908, f(x) = 0.6286
      10'h25E: recip_out = 32'h50698A86; // x = 0.5918, f(x) = 0.6282
      10'h25F: recip_out = 32'h505CEB70; // x = 0.5928, f(x) = 0.6278
      10'h260: recip_out = 32'h50505050; // x = 0.5938, f(x) = 0.6275
      10'h261: recip_out = 32'h5043B924; // x = 0.5947, f(x) = 0.6271
      10'h262: recip_out = 32'h503725EA; // x = 0.5957, f(x) = 0.6267
      10'h263: recip_out = 32'h502A96A0; // x = 0.5967, f(x) = 0.6263
      10'h264: recip_out = 32'h501E0B44; // x = 0.5977, f(x) = 0.6259
      10'h265: recip_out = 32'h501183D5; // x = 0.5986, f(x) = 0.6255
      10'h266: recip_out = 32'h50050050; // x = 0.5996, f(x) = 0.6252
      10'h267: recip_out = 32'h4FF880B4; // x = 0.6006, f(x) = 0.6248
      10'h268: recip_out = 32'h4FEC04FF; // x = 0.6016, f(x) = 0.6244
      10'h269: recip_out = 32'h4FDF8D2F; // x = 0.6025, f(x) = 0.6240
      10'h26A: recip_out = 32'h4FD31942; // x = 0.6035, f(x) = 0.6236
      10'h26B: recip_out = 32'h4FC6A936; // x = 0.6045, f(x) = 0.6233
      10'h26C: recip_out = 32'h4FBA3D0B; // x = 0.6055, f(x) = 0.6229
      10'h26D: recip_out = 32'h4FADD4BD; // x = 0.6064, f(x) = 0.6225
      10'h26E: recip_out = 32'h4FA1704B; // x = 0.6074, f(x) = 0.6221
      10'h26F: recip_out = 32'h4F950FB3; // x = 0.6084, f(x) = 0.6217
      10'h270: recip_out = 32'h4F88B2F4; // x = 0.6094, f(x) = 0.6214
      10'h271: recip_out = 32'h4F7C5A0B; // x = 0.6104, f(x) = 0.6210
      10'h272: recip_out = 32'h4F7004F7; // x = 0.6113, f(x) = 0.6206
      10'h273: recip_out = 32'h4F63B3B6; // x = 0.6123, f(x) = 0.6202
      10'h274: recip_out = 32'h4F576647; // x = 0.6133, f(x) = 0.6199
      10'h275: recip_out = 32'h4F4B1CA7; // x = 0.6143, f(x) = 0.6195
      10'h276: recip_out = 32'h4F3ED6D4; // x = 0.6152, f(x) = 0.6191
      10'h277: recip_out = 32'h4F3294CE; // x = 0.6162, f(x) = 0.6187
      10'h278: recip_out = 32'h4F265692; // x = 0.6172, f(x) = 0.6184
      10'h279: recip_out = 32'h4F1A1C1E; // x = 0.6182, f(x) = 0.6180
      10'h27A: recip_out = 32'h4F0DE571; // x = 0.6191, f(x) = 0.6176
      10'h27B: recip_out = 32'h4F01B289; // x = 0.6201, f(x) = 0.6172
      10'h27C: recip_out = 32'h4EF58365; // x = 0.6211, f(x) = 0.6169
      10'h27D: recip_out = 32'h4EE95801; // x = 0.6221, f(x) = 0.6165
      10'h27E: recip_out = 32'h4EDD305E; // x = 0.6230, f(x) = 0.6161
      10'h27F: recip_out = 32'h4ED10C78; // x = 0.6240, f(x) = 0.6158
      10'h280: recip_out = 32'h4EC4EC4F; // x = 0.6250, f(x) = 0.6154
      10'h281: recip_out = 32'h4EB8CFE0; // x = 0.6260, f(x) = 0.6150
      10'h282: recip_out = 32'h4EACB72A; // x = 0.6270, f(x) = 0.6146
      10'h283: recip_out = 32'h4EA0A22B; // x = 0.6279, f(x) = 0.6143
      10'h284: recip_out = 32'h4E9490E2; // x = 0.6289, f(x) = 0.6139
      10'h285: recip_out = 32'h4E88834C; // x = 0.6299, f(x) = 0.6135
      10'h286: recip_out = 32'h4E7C7969; // x = 0.6309, f(x) = 0.6132
      10'h287: recip_out = 32'h4E707335; // x = 0.6318, f(x) = 0.6128
      10'h288: recip_out = 32'h4E6470B0; // x = 0.6328, f(x) = 0.6124
      10'h289: recip_out = 32'h4E5871D9; // x = 0.6338, f(x) = 0.6121
      10'h28A: recip_out = 32'h4E4C76AC; // x = 0.6348, f(x) = 0.6117
      10'h28B: recip_out = 32'h4E407F29; // x = 0.6357, f(x) = 0.6113
      10'h28C: recip_out = 32'h4E348B4E; // x = 0.6367, f(x) = 0.6110
      10'h28D: recip_out = 32'h4E289B19; // x = 0.6377, f(x) = 0.6106
      10'h28E: recip_out = 32'h4E1CAE88; // x = 0.6387, f(x) = 0.6103
      10'h28F: recip_out = 32'h4E10C59A; // x = 0.6396, f(x) = 0.6099
      10'h290: recip_out = 32'h4E04E04E; // x = 0.6406, f(x) = 0.6095
      10'h291: recip_out = 32'h4DF8FEA1; // x = 0.6416, f(x) = 0.6092
      10'h292: recip_out = 32'h4DED2092; // x = 0.6426, f(x) = 0.6088
      10'h293: recip_out = 32'h4DE1461F; // x = 0.6436, f(x) = 0.6084
      10'h294: recip_out = 32'h4DD56F47; // x = 0.6445, f(x) = 0.6081
      10'h295: recip_out = 32'h4DC99C08; // x = 0.6455, f(x) = 0.6077
      10'h296: recip_out = 32'h4DBDCC60; // x = 0.6465, f(x) = 0.6074
      10'h297: recip_out = 32'h4DB2004E; // x = 0.6475, f(x) = 0.6070
      10'h298: recip_out = 32'h4DA637CF; // x = 0.6484, f(x) = 0.6066
      10'h299: recip_out = 32'h4D9A72E4; // x = 0.6494, f(x) = 0.6063
      10'h29A: recip_out = 32'h4D8EB189; // x = 0.6504, f(x) = 0.6059
      10'h29B: recip_out = 32'h4D82F3BD; // x = 0.6514, f(x) = 0.6056
      10'h29C: recip_out = 32'h4D77397E; // x = 0.6523, f(x) = 0.6052
      10'h29D: recip_out = 32'h4D6B82CC; // x = 0.6533, f(x) = 0.6048
      10'h29E: recip_out = 32'h4D5FCFA4; // x = 0.6543, f(x) = 0.6045
      10'h29F: recip_out = 32'h4D542005; // x = 0.6553, f(x) = 0.6041
      10'h2A0: recip_out = 32'h4D4873ED; // x = 0.6562, f(x) = 0.6038
      10'h2A1: recip_out = 32'h4D3CCB5A; // x = 0.6572, f(x) = 0.6034
      10'h2A2: recip_out = 32'h4D31264B; // x = 0.6582, f(x) = 0.6031
      10'h2A3: recip_out = 32'h4D2584BF; // x = 0.6592, f(x) = 0.6027
      10'h2A4: recip_out = 32'h4D19E6B4; // x = 0.6602, f(x) = 0.6024
      10'h2A5: recip_out = 32'h4D0E4C27; // x = 0.6611, f(x) = 0.6020
      10'h2A6: recip_out = 32'h4D02B518; // x = 0.6621, f(x) = 0.6016
      10'h2A7: recip_out = 32'h4CF72186; // x = 0.6631, f(x) = 0.6013
      10'h2A8: recip_out = 32'h4CEB916D; // x = 0.6641, f(x) = 0.6009
      10'h2A9: recip_out = 32'h4CE004CE; // x = 0.6650, f(x) = 0.6006
      10'h2AA: recip_out = 32'h4CD47BA6; // x = 0.6660, f(x) = 0.6002
      10'h2AB: recip_out = 32'h4CC8F5F4; // x = 0.6670, f(x) = 0.5999
      10'h2AC: recip_out = 32'h4CBD73B6; // x = 0.6680, f(x) = 0.5995
      10'h2AD: recip_out = 32'h4CB1F4EA; // x = 0.6689, f(x) = 0.5992
      10'h2AE: recip_out = 32'h4CA67990; // x = 0.6699, f(x) = 0.5988
      10'h2AF: recip_out = 32'h4C9B01A5; // x = 0.6709, f(x) = 0.5985
      10'h2B0: recip_out = 32'h4C8F8D29; // x = 0.6719, f(x) = 0.5981
      10'h2B1: recip_out = 32'h4C841C19; // x = 0.6729, f(x) = 0.5978
      10'h2B2: recip_out = 32'h4C78AE73; // x = 0.6738, f(x) = 0.5974
      10'h2B3: recip_out = 32'h4C6D4438; // x = 0.6748, f(x) = 0.5971
      10'h2B4: recip_out = 32'h4C61DD64; // x = 0.6758, f(x) = 0.5967
      10'h2B5: recip_out = 32'h4C5679F6; // x = 0.6768, f(x) = 0.5964
      10'h2B6: recip_out = 32'h4C4B19EE; // x = 0.6777, f(x) = 0.5960
      10'h2B7: recip_out = 32'h4C3FBD48; // x = 0.6787, f(x) = 0.5957
      10'h2B8: recip_out = 32'h4C346405; // x = 0.6797, f(x) = 0.5953
      10'h2B9: recip_out = 32'h4C290E22; // x = 0.6807, f(x) = 0.5950
      10'h2BA: recip_out = 32'h4C1DBB9D; // x = 0.6816, f(x) = 0.5947
      10'h2BB: recip_out = 32'h4C126C76; // x = 0.6826, f(x) = 0.5943
      10'h2BC: recip_out = 32'h4C0720AB; // x = 0.6836, f(x) = 0.5940
      10'h2BD: recip_out = 32'h4BFBD83A; // x = 0.6846, f(x) = 0.5936
      10'h2BE: recip_out = 32'h4BF09322; // x = 0.6855, f(x) = 0.5933
      10'h2BF: recip_out = 32'h4BE55161; // x = 0.6865, f(x) = 0.5929
      10'h2C0: recip_out = 32'h4BDA12F7; // x = 0.6875, f(x) = 0.5926
      10'h2C1: recip_out = 32'h4BCED7E0; // x = 0.6885, f(x) = 0.5922
      10'h2C2: recip_out = 32'h4BC3A01C; // x = 0.6895, f(x) = 0.5919
      10'h2C3: recip_out = 32'h4BB86BAA; // x = 0.6904, f(x) = 0.5916
      10'h2C4: recip_out = 32'h4BAD3A88; // x = 0.6914, f(x) = 0.5912
      10'h2C5: recip_out = 32'h4BA20CB4; // x = 0.6924, f(x) = 0.5909
      10'h2C6: recip_out = 32'h4B96E22D; // x = 0.6934, f(x) = 0.5905
      10'h2C7: recip_out = 32'h4B8BBAF2; // x = 0.6943, f(x) = 0.5902
      10'h2C8: recip_out = 32'h4B809701; // x = 0.6953, f(x) = 0.5899
      10'h2C9: recip_out = 32'h4B757659; // x = 0.6963, f(x) = 0.5895
      10'h2CA: recip_out = 32'h4B6A58F7; // x = 0.6973, f(x) = 0.5892
      10'h2CB: recip_out = 32'h4B5F3EDC; // x = 0.6982, f(x) = 0.5888
      10'h2CC: recip_out = 32'h4B542805; // x = 0.6992, f(x) = 0.5885
      10'h2CD: recip_out = 32'h4B491470; // x = 0.7002, f(x) = 0.5882
      10'h2CE: recip_out = 32'h4B3E041D; // x = 0.7012, f(x) = 0.5878
      10'h2CF: recip_out = 32'h4B32F70A; // x = 0.7021, f(x) = 0.5875
      10'h2D0: recip_out = 32'h4B27ED36; // x = 0.7031, f(x) = 0.5872
      10'h2D1: recip_out = 32'h4B1CE69F; // x = 0.7041, f(x) = 0.5868
      10'h2D2: recip_out = 32'h4B11E343; // x = 0.7051, f(x) = 0.5865
      10'h2D3: recip_out = 32'h4B06E322; // x = 0.7061, f(x) = 0.5861
      10'h2D4: recip_out = 32'h4AFBE639; // x = 0.7070, f(x) = 0.5858
      10'h2D5: recip_out = 32'h4AF0EC88; // x = 0.7080, f(x) = 0.5855
      10'h2D6: recip_out = 32'h4AE5F60D; // x = 0.7090, f(x) = 0.5851
      10'h2D7: recip_out = 32'h4ADB02C7; // x = 0.7100, f(x) = 0.5848
      10'h2D8: recip_out = 32'h4AD012B4; // x = 0.7109, f(x) = 0.5845
      10'h2D9: recip_out = 32'h4AC525D3; // x = 0.7119, f(x) = 0.5841
      10'h2DA: recip_out = 32'h4ABA3C22; // x = 0.7129, f(x) = 0.5838
      10'h2DB: recip_out = 32'h4AAF55A0; // x = 0.7139, f(x) = 0.5835
      10'h2DC: recip_out = 32'h4AA4724C; // x = 0.7148, f(x) = 0.5831
      10'h2DD: recip_out = 32'h4A999224; // x = 0.7158, f(x) = 0.5828
      10'h2DE: recip_out = 32'h4A8EB527; // x = 0.7168, f(x) = 0.5825
      10'h2DF: recip_out = 32'h4A83DB53; // x = 0.7178, f(x) = 0.5821
      10'h2E0: recip_out = 32'h4A7904A8; // x = 0.7188, f(x) = 0.5818
      10'h2E1: recip_out = 32'h4A6E3123; // x = 0.7197, f(x) = 0.5815
      10'h2E2: recip_out = 32'h4A6360C3; // x = 0.7207, f(x) = 0.5812
      10'h2E3: recip_out = 32'h4A589388; // x = 0.7217, f(x) = 0.5808
      10'h2E4: recip_out = 32'h4A4DC96F; // x = 0.7227, f(x) = 0.5805
      10'h2E5: recip_out = 32'h4A430277; // x = 0.7236, f(x) = 0.5802
      10'h2E6: recip_out = 32'h4A383E9F; // x = 0.7246, f(x) = 0.5798
      10'h2E7: recip_out = 32'h4A2D7DE6; // x = 0.7256, f(x) = 0.5795
      10'h2E8: recip_out = 32'h4A22C04A; // x = 0.7266, f(x) = 0.5792
      10'h2E9: recip_out = 32'h4A1805CA; // x = 0.7275, f(x) = 0.5789
      10'h2EA: recip_out = 32'h4A0D4E64; // x = 0.7285, f(x) = 0.5785
      10'h2EB: recip_out = 32'h4A029A17; // x = 0.7295, f(x) = 0.5782
      10'h2EC: recip_out = 32'h49F7E8E3; // x = 0.7305, f(x) = 0.5779
      10'h2ED: recip_out = 32'h49ED3AC4; // x = 0.7314, f(x) = 0.5776
      10'h2EE: recip_out = 32'h49E28FBB; // x = 0.7324, f(x) = 0.5772
      10'h2EF: recip_out = 32'h49D7E7C5; // x = 0.7334, f(x) = 0.5769
      10'h2F0: recip_out = 32'h49CD42E2; // x = 0.7344, f(x) = 0.5766
      10'h2F1: recip_out = 32'h49C2A110; // x = 0.7354, f(x) = 0.5763
      10'h2F2: recip_out = 32'h49B8024E; // x = 0.7363, f(x) = 0.5759
      10'h2F3: recip_out = 32'h49AD669A; // x = 0.7373, f(x) = 0.5756
      10'h2F4: recip_out = 32'h49A2CDF3; // x = 0.7383, f(x) = 0.5753
      10'h2F5: recip_out = 32'h49983859; // x = 0.7393, f(x) = 0.5750
      10'h2F6: recip_out = 32'h498DA5C8; // x = 0.7402, f(x) = 0.5746
      10'h2F7: recip_out = 32'h49831641; // x = 0.7412, f(x) = 0.5743
      10'h2F8: recip_out = 32'h497889C2; // x = 0.7422, f(x) = 0.5740
      10'h2F9: recip_out = 32'h496E0049; // x = 0.7432, f(x) = 0.5737
      10'h2FA: recip_out = 32'h496379D6; // x = 0.7441, f(x) = 0.5733
      10'h2FB: recip_out = 32'h4958F667; // x = 0.7451, f(x) = 0.5730
      10'h2FC: recip_out = 32'h494E75FA; // x = 0.7461, f(x) = 0.5727
      10'h2FD: recip_out = 32'h4943F88F; // x = 0.7471, f(x) = 0.5724
      10'h2FE: recip_out = 32'h49397E24; // x = 0.7480, f(x) = 0.5721
      10'h2FF: recip_out = 32'h492F06B8; // x = 0.7490, f(x) = 0.5717
      10'h300: recip_out = 32'h49249249; // x = 0.7500, f(x) = 0.5714
      10'h301: recip_out = 32'h491A20D7; // x = 0.7510, f(x) = 0.5711
      10'h302: recip_out = 32'h490FB25F; // x = 0.7520, f(x) = 0.5708
      10'h303: recip_out = 32'h490546E2; // x = 0.7529, f(x) = 0.5705
      10'h304: recip_out = 32'h48FADE5C; // x = 0.7539, f(x) = 0.5702
      10'h305: recip_out = 32'h48F078CE; // x = 0.7549, f(x) = 0.5698
      10'h306: recip_out = 32'h48E61636; // x = 0.7559, f(x) = 0.5695
      10'h307: recip_out = 32'h48DBB693; // x = 0.7568, f(x) = 0.5692
      10'h308: recip_out = 32'h48D159E2; // x = 0.7578, f(x) = 0.5689
      10'h309: recip_out = 32'h48C70024; // x = 0.7588, f(x) = 0.5686
      10'h30A: recip_out = 32'h48BCA957; // x = 0.7598, f(x) = 0.5683
      10'h30B: recip_out = 32'h48B2557A; // x = 0.7607, f(x) = 0.5679
      10'h30C: recip_out = 32'h48A8048B; // x = 0.7617, f(x) = 0.5676
      10'h30D: recip_out = 32'h489DB688; // x = 0.7627, f(x) = 0.5673
      10'h30E: recip_out = 32'h48936B72; // x = 0.7637, f(x) = 0.5670
      10'h30F: recip_out = 32'h48892347; // x = 0.7646, f(x) = 0.5667
      10'h310: recip_out = 32'h487EDE05; // x = 0.7656, f(x) = 0.5664
      10'h311: recip_out = 32'h48749BAB; // x = 0.7666, f(x) = 0.5661
      10'h312: recip_out = 32'h486A5C37; // x = 0.7676, f(x) = 0.5657
      10'h313: recip_out = 32'h48601FAA; // x = 0.7686, f(x) = 0.5654
      10'h314: recip_out = 32'h4855E601; // x = 0.7695, f(x) = 0.5651
      10'h315: recip_out = 32'h484BAF3B; // x = 0.7705, f(x) = 0.5648
      10'h316: recip_out = 32'h48417B58; // x = 0.7715, f(x) = 0.5645
      10'h317: recip_out = 32'h48374A55; // x = 0.7725, f(x) = 0.5642
      10'h318: recip_out = 32'h482D1C32; // x = 0.7734, f(x) = 0.5639
      10'h319: recip_out = 32'h4822F0ED; // x = 0.7744, f(x) = 0.5636
      10'h31A: recip_out = 32'h4818C885; // x = 0.7754, f(x) = 0.5633
      10'h31B: recip_out = 32'h480EA2F9; // x = 0.7764, f(x) = 0.5629
      10'h31C: recip_out = 32'h48048048; // x = 0.7773, f(x) = 0.5626
      10'h31D: recip_out = 32'h47FA6070; // x = 0.7783, f(x) = 0.5623
      10'h31E: recip_out = 32'h47F04371; // x = 0.7793, f(x) = 0.5620
      10'h31F: recip_out = 32'h47E62949; // x = 0.7803, f(x) = 0.5617
      10'h320: recip_out = 32'h47DC11F7; // x = 0.7812, f(x) = 0.5614
      10'h321: recip_out = 32'h47D1FD7A; // x = 0.7822, f(x) = 0.5611
      10'h322: recip_out = 32'h47C7EBD0; // x = 0.7832, f(x) = 0.5608
      10'h323: recip_out = 32'h47BDDCF8; // x = 0.7842, f(x) = 0.5605
      10'h324: recip_out = 32'h47B3D0F2; // x = 0.7852, f(x) = 0.5602
      10'h325: recip_out = 32'h47A9C7BC; // x = 0.7861, f(x) = 0.5599
      10'h326: recip_out = 32'h479FC154; // x = 0.7871, f(x) = 0.5596
      10'h327: recip_out = 32'h4795BDBA; // x = 0.7881, f(x) = 0.5593
      10'h328: recip_out = 32'h478BBCED; // x = 0.7891, f(x) = 0.5590
      10'h329: recip_out = 32'h4781BEEB; // x = 0.7900, f(x) = 0.5586
      10'h32A: recip_out = 32'h4777C3B3; // x = 0.7910, f(x) = 0.5583
      10'h32B: recip_out = 32'h476DCB44; // x = 0.7920, f(x) = 0.5580
      10'h32C: recip_out = 32'h4763D59D; // x = 0.7930, f(x) = 0.5577
      10'h32D: recip_out = 32'h4759E2BC; // x = 0.7939, f(x) = 0.5574
      10'h32E: recip_out = 32'h474FF2A1; // x = 0.7949, f(x) = 0.5571
      10'h32F: recip_out = 32'h4746054A; // x = 0.7959, f(x) = 0.5568
      10'h330: recip_out = 32'h473C1AB7; // x = 0.7969, f(x) = 0.5565
      10'h331: recip_out = 32'h473232E5; // x = 0.7979, f(x) = 0.5562
      10'h332: recip_out = 32'h47284DD4; // x = 0.7988, f(x) = 0.5559
      10'h333: recip_out = 32'h471E6B83; // x = 0.7998, f(x) = 0.5556
      10'h334: recip_out = 32'h47148BF0; // x = 0.8008, f(x) = 0.5553
      10'h335: recip_out = 32'h470AAF1B; // x = 0.8018, f(x) = 0.5550
      10'h336: recip_out = 32'h4700D502; // x = 0.8027, f(x) = 0.5547
      10'h337: recip_out = 32'h46F6FDA5; // x = 0.8037, f(x) = 0.5544
      10'h338: recip_out = 32'h46ED2901; // x = 0.8047, f(x) = 0.5541
      10'h339: recip_out = 32'h46E35716; // x = 0.8057, f(x) = 0.5538
      10'h33A: recip_out = 32'h46D987E3; // x = 0.8066, f(x) = 0.5535
      10'h33B: recip_out = 32'h46CFBB67; // x = 0.8076, f(x) = 0.5532
      10'h33C: recip_out = 32'h46C5F1A0; // x = 0.8086, f(x) = 0.5529
      10'h33D: recip_out = 32'h46BC2A8D; // x = 0.8096, f(x) = 0.5526
      10'h33E: recip_out = 32'h46B2662E; // x = 0.8105, f(x) = 0.5523
      10'h33F: recip_out = 32'h46A8A481; // x = 0.8115, f(x) = 0.5520
      10'h340: recip_out = 32'h469EE584; // x = 0.8125, f(x) = 0.5517
      10'h341: recip_out = 32'h46952938; // x = 0.8135, f(x) = 0.5514
      10'h342: recip_out = 32'h468B6F9B; // x = 0.8145, f(x) = 0.5511
      10'h343: recip_out = 32'h4681B8AB; // x = 0.8154, f(x) = 0.5508
      10'h344: recip_out = 32'h46780468; // x = 0.8164, f(x) = 0.5505
      10'h345: recip_out = 32'h466E52D0; // x = 0.8174, f(x) = 0.5502
      10'h346: recip_out = 32'h4664A3E2; // x = 0.8184, f(x) = 0.5499
      10'h347: recip_out = 32'h465AF79E; // x = 0.8193, f(x) = 0.5497
      10'h348: recip_out = 32'h46514E02; // x = 0.8203, f(x) = 0.5494
      10'h349: recip_out = 32'h4647A70D; // x = 0.8213, f(x) = 0.5491
      10'h34A: recip_out = 32'h463E02BE; // x = 0.8223, f(x) = 0.5488
      10'h34B: recip_out = 32'h46346114; // x = 0.8232, f(x) = 0.5485
      10'h34C: recip_out = 32'h462AC20E; // x = 0.8242, f(x) = 0.5482
      10'h34D: recip_out = 32'h462125AB; // x = 0.8252, f(x) = 0.5479
      10'h34E: recip_out = 32'h46178BE9; // x = 0.8262, f(x) = 0.5476
      10'h34F: recip_out = 32'h460DF4C8; // x = 0.8271, f(x) = 0.5473
      10'h350: recip_out = 32'h46046046; // x = 0.8281, f(x) = 0.5470
      10'h351: recip_out = 32'h45FACE63; // x = 0.8291, f(x) = 0.5467
      10'h352: recip_out = 32'h45F13F1D; // x = 0.8301, f(x) = 0.5464
      10'h353: recip_out = 32'h45E7B273; // x = 0.8311, f(x) = 0.5461
      10'h354: recip_out = 32'h45DE2864; // x = 0.8320, f(x) = 0.5458
      10'h355: recip_out = 32'h45D4A0F0; // x = 0.8330, f(x) = 0.5456
      10'h356: recip_out = 32'h45CB1C15; // x = 0.8340, f(x) = 0.5453
      10'h357: recip_out = 32'h45C199D1; // x = 0.8350, f(x) = 0.5450
      10'h358: recip_out = 32'h45B81A25; // x = 0.8359, f(x) = 0.5447
      10'h359: recip_out = 32'h45AE9D0F; // x = 0.8369, f(x) = 0.5444
      10'h35A: recip_out = 32'h45A5228D; // x = 0.8379, f(x) = 0.5441
      10'h35B: recip_out = 32'h459BAA9F; // x = 0.8389, f(x) = 0.5438
      10'h35C: recip_out = 32'h45923544; // x = 0.8398, f(x) = 0.5435
      10'h35D: recip_out = 32'h4588C27A; // x = 0.8408, f(x) = 0.5432
      10'h35E: recip_out = 32'h457F5242; // x = 0.8418, f(x) = 0.5429
      10'h35F: recip_out = 32'h4575E498; // x = 0.8428, f(x) = 0.5427
      10'h360: recip_out = 32'h456C797E; // x = 0.8438, f(x) = 0.5424
      10'h361: recip_out = 32'h456310F1; // x = 0.8447, f(x) = 0.5421
      10'h362: recip_out = 32'h4559AAF0; // x = 0.8457, f(x) = 0.5418
      10'h363: recip_out = 32'h4550477B; // x = 0.8467, f(x) = 0.5415
      10'h364: recip_out = 32'h4546E690; // x = 0.8477, f(x) = 0.5412
      10'h365: recip_out = 32'h453D882F; // x = 0.8486, f(x) = 0.5409
      10'h366: recip_out = 32'h45342C55; // x = 0.8496, f(x) = 0.5407
      10'h367: recip_out = 32'h452AD304; // x = 0.8506, f(x) = 0.5404
      10'h368: recip_out = 32'h45217C38; // x = 0.8516, f(x) = 0.5401
      10'h369: recip_out = 32'h451827F2; // x = 0.8525, f(x) = 0.5398
      10'h36A: recip_out = 32'h450ED630; // x = 0.8535, f(x) = 0.5395
      10'h36B: recip_out = 32'h450586F1; // x = 0.8545, f(x) = 0.5392
      10'h36C: recip_out = 32'h44FC3A35; // x = 0.8555, f(x) = 0.5389
      10'h36D: recip_out = 32'h44F2EFFA; // x = 0.8564, f(x) = 0.5387
      10'h36E: recip_out = 32'h44E9A83E; // x = 0.8574, f(x) = 0.5384
      10'h36F: recip_out = 32'h44E06303; // x = 0.8584, f(x) = 0.5381
      10'h370: recip_out = 32'h44D72045; // x = 0.8594, f(x) = 0.5378
      10'h371: recip_out = 32'h44CDE004; // x = 0.8604, f(x) = 0.5375
      10'h372: recip_out = 32'h44C4A240; // x = 0.8613, f(x) = 0.5373
      10'h373: recip_out = 32'h44BB66F7; // x = 0.8623, f(x) = 0.5370
      10'h374: recip_out = 32'h44B22E28; // x = 0.8633, f(x) = 0.5367
      10'h375: recip_out = 32'h44A8F7D2; // x = 0.8643, f(x) = 0.5364
      10'h376: recip_out = 32'h449FC3F4; // x = 0.8652, f(x) = 0.5361
      10'h377: recip_out = 32'h4496928E; // x = 0.8662, f(x) = 0.5358
      10'h378: recip_out = 32'h448D639D; // x = 0.8672, f(x) = 0.5356
      10'h379: recip_out = 32'h44843722; // x = 0.8682, f(x) = 0.5353
      10'h37A: recip_out = 32'h447B0D1C; // x = 0.8691, f(x) = 0.5350
      10'h37B: recip_out = 32'h4471E588; // x = 0.8701, f(x) = 0.5347
      10'h37C: recip_out = 32'h4468C067; // x = 0.8711, f(x) = 0.5344
      10'h37D: recip_out = 32'h445F9DB7; // x = 0.8721, f(x) = 0.5342
      10'h37E: recip_out = 32'h44567D77; // x = 0.8730, f(x) = 0.5339
      10'h37F: recip_out = 32'h444D5FA6; // x = 0.8740, f(x) = 0.5336
      10'h380: recip_out = 32'h44444444; // x = 0.8750, f(x) = 0.5333
      10'h381: recip_out = 32'h443B2B50; // x = 0.8760, f(x) = 0.5331
      10'h382: recip_out = 32'h443214C7; // x = 0.8770, f(x) = 0.5328
      10'h383: recip_out = 32'h442900AA; // x = 0.8779, f(x) = 0.5325
      10'h384: recip_out = 32'h441FEEF8; // x = 0.8789, f(x) = 0.5322
      10'h385: recip_out = 32'h4416DFAF; // x = 0.8799, f(x) = 0.5319
      10'h386: recip_out = 32'h440DD2CF; // x = 0.8809, f(x) = 0.5317
      10'h387: recip_out = 32'h4404C856; // x = 0.8818, f(x) = 0.5314
      10'h388: recip_out = 32'h43FBC044; // x = 0.8828, f(x) = 0.5311
      10'h389: recip_out = 32'h43F2BA98; // x = 0.8838, f(x) = 0.5308
      10'h38A: recip_out = 32'h43E9B750; // x = 0.8848, f(x) = 0.5306
      10'h38B: recip_out = 32'h43E0B66C; // x = 0.8857, f(x) = 0.5303
      10'h38C: recip_out = 32'h43D7B7EB; // x = 0.8867, f(x) = 0.5300
      10'h38D: recip_out = 32'h43CEBBCC; // x = 0.8877, f(x) = 0.5297
      10'h38E: recip_out = 32'h43C5C20D; // x = 0.8887, f(x) = 0.5295
      10'h38F: recip_out = 32'h43BCCAAF; // x = 0.8896, f(x) = 0.5292
      10'h390: recip_out = 32'h43B3D5B0; // x = 0.8906, f(x) = 0.5289
      10'h391: recip_out = 32'h43AAE30E; // x = 0.8916, f(x) = 0.5287
      10'h392: recip_out = 32'h43A1F2CA; // x = 0.8926, f(x) = 0.5284
      10'h393: recip_out = 32'h439904E3; // x = 0.8936, f(x) = 0.5281
      10'h394: recip_out = 32'h43901956; // x = 0.8945, f(x) = 0.5278
      10'h395: recip_out = 32'h43873024; // x = 0.8955, f(x) = 0.5276
      10'h396: recip_out = 32'h437E494B; // x = 0.8965, f(x) = 0.5273
      10'h397: recip_out = 32'h437564CB; // x = 0.8975, f(x) = 0.5270
      10'h398: recip_out = 32'h436C82A2; // x = 0.8984, f(x) = 0.5267
      10'h399: recip_out = 32'h4363A2D0; // x = 0.8994, f(x) = 0.5265
      10'h39A: recip_out = 32'h435AC554; // x = 0.9004, f(x) = 0.5262
      10'h39B: recip_out = 32'h4351EA2C; // x = 0.9014, f(x) = 0.5259
      10'h39C: recip_out = 32'h43491159; // x = 0.9023, f(x) = 0.5257
      10'h39D: recip_out = 32'h43403AD8; // x = 0.9033, f(x) = 0.5254
      10'h39E: recip_out = 32'h433766AA; // x = 0.9043, f(x) = 0.5251
      10'h39F: recip_out = 32'h432E94CC; // x = 0.9053, f(x) = 0.5249
      10'h3A0: recip_out = 32'h4325C53F; // x = 0.9062, f(x) = 0.5246
      10'h3A1: recip_out = 32'h431CF801; // x = 0.9072, f(x) = 0.5243
      10'h3A2: recip_out = 32'h43142D12; // x = 0.9082, f(x) = 0.5241
      10'h3A3: recip_out = 32'h430B6470; // x = 0.9092, f(x) = 0.5238
      10'h3A4: recip_out = 32'h43029E1A; // x = 0.9102, f(x) = 0.5235
      10'h3A5: recip_out = 32'h42F9DA10; // x = 0.9111, f(x) = 0.5232
      10'h3A6: recip_out = 32'h42F11852; // x = 0.9121, f(x) = 0.5230
      10'h3A7: recip_out = 32'h42E858DD; // x = 0.9131, f(x) = 0.5227
      10'h3A8: recip_out = 32'h42DF9BB1; // x = 0.9141, f(x) = 0.5224
      10'h3A9: recip_out = 32'h42D6E0CD; // x = 0.9150, f(x) = 0.5222
      10'h3AA: recip_out = 32'h42CE2830; // x = 0.9160, f(x) = 0.5219
      10'h3AB: recip_out = 32'h42C571DA; // x = 0.9170, f(x) = 0.5217
      10'h3AC: recip_out = 32'h42BCBDC9; // x = 0.9180, f(x) = 0.5214
      10'h3AD: recip_out = 32'h42B40BFC; // x = 0.9189, f(x) = 0.5211
      10'h3AE: recip_out = 32'h42AB5C74; // x = 0.9199, f(x) = 0.5209
      10'h3AF: recip_out = 32'h42A2AF2E; // x = 0.9209, f(x) = 0.5206
      10'h3B0: recip_out = 32'h429A042A; // x = 0.9219, f(x) = 0.5203
      10'h3B1: recip_out = 32'h42915B67; // x = 0.9229, f(x) = 0.5201
      10'h3B2: recip_out = 32'h4288B4E4; // x = 0.9238, f(x) = 0.5198
      10'h3B3: recip_out = 32'h428010A0; // x = 0.9248, f(x) = 0.5195
      10'h3B4: recip_out = 32'h42776E9B; // x = 0.9258, f(x) = 0.5193
      10'h3B5: recip_out = 32'h426ECED3; // x = 0.9268, f(x) = 0.5190
      10'h3B6: recip_out = 32'h42663148; // x = 0.9277, f(x) = 0.5187
      10'h3B7: recip_out = 32'h425D95F8; // x = 0.9287, f(x) = 0.5185
      10'h3B8: recip_out = 32'h4254FCE4; // x = 0.9297, f(x) = 0.5182
      10'h3B9: recip_out = 32'h424C660A; // x = 0.9307, f(x) = 0.5180
      10'h3BA: recip_out = 32'h4243D168; // x = 0.9316, f(x) = 0.5177
      10'h3BB: recip_out = 32'h423B3EFF; // x = 0.9326, f(x) = 0.5174
      10'h3BC: recip_out = 32'h4232AECE; // x = 0.9336, f(x) = 0.5172
      10'h3BD: recip_out = 32'h422A20D3; // x = 0.9346, f(x) = 0.5169
      10'h3BE: recip_out = 32'h4221950E; // x = 0.9355, f(x) = 0.5166
      10'h3BF: recip_out = 32'h42190B7D; // x = 0.9365, f(x) = 0.5164
      10'h3C0: recip_out = 32'h42108421; // x = 0.9375, f(x) = 0.5161
      10'h3C1: recip_out = 32'h4207FEF8; // x = 0.9385, f(x) = 0.5159
      10'h3C2: recip_out = 32'h41FF7C01; // x = 0.9395, f(x) = 0.5156
      10'h3C3: recip_out = 32'h41F6FB3C; // x = 0.9404, f(x) = 0.5153
      10'h3C4: recip_out = 32'h41EE7CA7; // x = 0.9414, f(x) = 0.5151
      10'h3C5: recip_out = 32'h41E60042; // x = 0.9424, f(x) = 0.5148
      10'h3C6: recip_out = 32'h41DD860C; // x = 0.9434, f(x) = 0.5146
      10'h3C7: recip_out = 32'h41D50E04; // x = 0.9443, f(x) = 0.5143
      10'h3C8: recip_out = 32'h41CC9829; // x = 0.9453, f(x) = 0.5141
      10'h3C9: recip_out = 32'h41C4247B; // x = 0.9463, f(x) = 0.5138
      10'h3CA: recip_out = 32'h41BBB2F8; // x = 0.9473, f(x) = 0.5135
      10'h3CB: recip_out = 32'h41B343A0; // x = 0.9482, f(x) = 0.5133
      10'h3CC: recip_out = 32'h41AAD672; // x = 0.9492, f(x) = 0.5130
      10'h3CD: recip_out = 32'h41A26B6D; // x = 0.9502, f(x) = 0.5128
      10'h3CE: recip_out = 32'h419A0290; // x = 0.9512, f(x) = 0.5125
      10'h3CF: recip_out = 32'h41919BDB; // x = 0.9521, f(x) = 0.5123
      10'h3D0: recip_out = 32'h4189374C; // x = 0.9531, f(x) = 0.5120
      10'h3D1: recip_out = 32'h4180D4E3; // x = 0.9541, f(x) = 0.5117
      10'h3D2: recip_out = 32'h4178749F; // x = 0.9551, f(x) = 0.5115
      10'h3D3: recip_out = 32'h4170167F; // x = 0.9561, f(x) = 0.5112
      10'h3D4: recip_out = 32'h4167BA82; // x = 0.9570, f(x) = 0.5110
      10'h3D5: recip_out = 32'h415F60A8; // x = 0.9580, f(x) = 0.5107
      10'h3D6: recip_out = 32'h415708EF; // x = 0.9590, f(x) = 0.5105
      10'h3D7: recip_out = 32'h414EB357; // x = 0.9600, f(x) = 0.5102
      10'h3D8: recip_out = 32'h41465FDF; // x = 0.9609, f(x) = 0.5100
      10'h3D9: recip_out = 32'h413E0E87; // x = 0.9619, f(x) = 0.5097
      10'h3DA: recip_out = 32'h4135BF4D; // x = 0.9629, f(x) = 0.5095
      10'h3DB: recip_out = 32'h412D7230; // x = 0.9639, f(x) = 0.5092
      10'h3DC: recip_out = 32'h41252730; // x = 0.9648, f(x) = 0.5089
      10'h3DD: recip_out = 32'h411CDE4D; // x = 0.9658, f(x) = 0.5087
      10'h3DE: recip_out = 32'h41149784; // x = 0.9668, f(x) = 0.5084
      10'h3DF: recip_out = 32'h410C52D6; // x = 0.9678, f(x) = 0.5082
      10'h3E0: recip_out = 32'h41041041; // x = 0.9688, f(x) = 0.5079
      10'h3E1: recip_out = 32'h40FBCFC5; // x = 0.9697, f(x) = 0.5077
      10'h3E2: recip_out = 32'h40F39161; // x = 0.9707, f(x) = 0.5074
      10'h3E3: recip_out = 32'h40EB5514; // x = 0.9717, f(x) = 0.5072
      10'h3E4: recip_out = 32'h40E31ADE; // x = 0.9727, f(x) = 0.5069
      10'h3E5: recip_out = 32'h40DAE2BD; // x = 0.9736, f(x) = 0.5067
      10'h3E6: recip_out = 32'h40D2ACB1; // x = 0.9746, f(x) = 0.5064
      10'h3E7: recip_out = 32'h40CA78B9; // x = 0.9756, f(x) = 0.5062
      10'h3E8: recip_out = 32'h40C246D4; // x = 0.9766, f(x) = 0.5059
      10'h3E9: recip_out = 32'h40BA1702; // x = 0.9775, f(x) = 0.5057
      10'h3EA: recip_out = 32'h40B1E941; // x = 0.9785, f(x) = 0.5054
      10'h3EB: recip_out = 32'h40A9BD92; // x = 0.9795, f(x) = 0.5052
      10'h3EC: recip_out = 32'h40A193F2; // x = 0.9805, f(x) = 0.5049
      10'h3ED: recip_out = 32'h40996C61; // x = 0.9814, f(x) = 0.5047
      10'h3EE: recip_out = 32'h409146DF; // x = 0.9824, f(x) = 0.5044
      10'h3EF: recip_out = 32'h4089236B; // x = 0.9834, f(x) = 0.5042
      10'h3F0: recip_out = 32'h40810204; // x = 0.9844, f(x) = 0.5039
      10'h3F1: recip_out = 32'h4078E2A9; // x = 0.9854, f(x) = 0.5037
      10'h3F2: recip_out = 32'h4070C559; // x = 0.9863, f(x) = 0.5034
      10'h3F3: recip_out = 32'h4068AA14; // x = 0.9873, f(x) = 0.5032
      10'h3F4: recip_out = 32'h406090D9; // x = 0.9883, f(x) = 0.5029
      10'h3F5: recip_out = 32'h405879A7; // x = 0.9893, f(x) = 0.5027
      10'h3F6: recip_out = 32'h4050647E; // x = 0.9902, f(x) = 0.5025
      10'h3F7: recip_out = 32'h4048515C; // x = 0.9912, f(x) = 0.5022
      10'h3F8: recip_out = 32'h40404040; // x = 0.9922, f(x) = 0.5020
      10'h3F9: recip_out = 32'h4038312B; // x = 0.9932, f(x) = 0.5017
      10'h3FA: recip_out = 32'h4030241B; // x = 0.9941, f(x) = 0.5015
      10'h3FB: recip_out = 32'h40281910; // x = 0.9951, f(x) = 0.5012
      10'h3FC: recip_out = 32'h40201008; // x = 0.9961, f(x) = 0.5010
      10'h3FD: recip_out = 32'h40180903; // x = 0.9971, f(x) = 0.5007
      10'h3FE: recip_out = 32'h40100401; // x = 0.9980, f(x) = 0.5005
      10'h3FF: recip_out = 32'h40080100; // x = 0.9990, f(x) = 0.5002
      default: recip_out = 32'h00000000;
    endcase
end


wire [11:0] exp_addr = input_data0[31:20];
reg  [31:0] exp_out;
always @( * ) begin
        case ( exp_addr )
          12'h000: exp_out = 32'h7FFFFFFF; 
          12'h800: exp_out = 32'h000000F2; // x = -16.0000, f(x) = 0.0000
          12'h801: exp_out = 32'h000000F4; // x = -15.9922, f(x) = 0.0000
          12'h802: exp_out = 32'h000000F5; // x = -15.9844, f(x) = 0.0000
          12'h803: exp_out = 32'h000000F7; // x = -15.9766, f(x) = 0.0000
          12'h804: exp_out = 32'h000000F9; // x = -15.9688, f(x) = 0.0000
          12'h805: exp_out = 32'h000000FB; // x = -15.9609, f(x) = 0.0000
          12'h806: exp_out = 32'h000000FD; // x = -15.9531, f(x) = 0.0000
          12'h807: exp_out = 32'h000000FF; // x = -15.9453, f(x) = 0.0000
          12'h808: exp_out = 32'h00000101; // x = -15.9375, f(x) = 0.0000
          12'h809: exp_out = 32'h00000103; // x = -15.9297, f(x) = 0.0000
          12'h80A: exp_out = 32'h00000105; // x = -15.9219, f(x) = 0.0000
          12'h80B: exp_out = 32'h00000107; // x = -15.9141, f(x) = 0.0000
          12'h80C: exp_out = 32'h00000109; // x = -15.9062, f(x) = 0.0000
          12'h80D: exp_out = 32'h0000010C; // x = -15.8984, f(x) = 0.0000
          12'h80E: exp_out = 32'h0000010E; // x = -15.8906, f(x) = 0.0000
          12'h80F: exp_out = 32'h00000110; // x = -15.8828, f(x) = 0.0000
          12'h810: exp_out = 32'h00000112; // x = -15.8750, f(x) = 0.0000
          12'h811: exp_out = 32'h00000114; // x = -15.8672, f(x) = 0.0000
          12'h812: exp_out = 32'h00000116; // x = -15.8594, f(x) = 0.0000
          12'h813: exp_out = 32'h00000118; // x = -15.8516, f(x) = 0.0000
          12'h814: exp_out = 32'h0000011B; // x = -15.8438, f(x) = 0.0000
          12'h815: exp_out = 32'h0000011D; // x = -15.8359, f(x) = 0.0000
          12'h816: exp_out = 32'h0000011F; // x = -15.8281, f(x) = 0.0000
          12'h817: exp_out = 32'h00000121; // x = -15.8203, f(x) = 0.0000
          12'h818: exp_out = 32'h00000124; // x = -15.8125, f(x) = 0.0000
          12'h819: exp_out = 32'h00000126; // x = -15.8047, f(x) = 0.0000
          12'h81A: exp_out = 32'h00000128; // x = -15.7969, f(x) = 0.0000
          12'h81B: exp_out = 32'h0000012A; // x = -15.7891, f(x) = 0.0000
          12'h81C: exp_out = 32'h0000012D; // x = -15.7812, f(x) = 0.0000
          12'h81D: exp_out = 32'h0000012F; // x = -15.7734, f(x) = 0.0000
          12'h81E: exp_out = 32'h00000131; // x = -15.7656, f(x) = 0.0000
          12'h81F: exp_out = 32'h00000134; // x = -15.7578, f(x) = 0.0000
          12'h820: exp_out = 32'h00000136; // x = -15.7500, f(x) = 0.0000
          12'h821: exp_out = 32'h00000139; // x = -15.7422, f(x) = 0.0000
          12'h822: exp_out = 32'h0000013B; // x = -15.7344, f(x) = 0.0000
          12'h823: exp_out = 32'h0000013E; // x = -15.7266, f(x) = 0.0000
          12'h824: exp_out = 32'h00000140; // x = -15.7188, f(x) = 0.0000
          12'h825: exp_out = 32'h00000143; // x = -15.7109, f(x) = 0.0000
          12'h826: exp_out = 32'h00000145; // x = -15.7031, f(x) = 0.0000
          12'h827: exp_out = 32'h00000148; // x = -15.6953, f(x) = 0.0000
          12'h828: exp_out = 32'h0000014A; // x = -15.6875, f(x) = 0.0000
          12'h829: exp_out = 32'h0000014D; // x = -15.6797, f(x) = 0.0000
          12'h82A: exp_out = 32'h00000150; // x = -15.6719, f(x) = 0.0000
          12'h82B: exp_out = 32'h00000152; // x = -15.6641, f(x) = 0.0000
          12'h82C: exp_out = 32'h00000155; // x = -15.6562, f(x) = 0.0000
          12'h82D: exp_out = 32'h00000157; // x = -15.6484, f(x) = 0.0000
          12'h82E: exp_out = 32'h0000015A; // x = -15.6406, f(x) = 0.0000
          12'h82F: exp_out = 32'h0000015D; // x = -15.6328, f(x) = 0.0000
          12'h830: exp_out = 32'h00000160; // x = -15.6250, f(x) = 0.0000
          12'h831: exp_out = 32'h00000162; // x = -15.6172, f(x) = 0.0000
          12'h832: exp_out = 32'h00000165; // x = -15.6094, f(x) = 0.0000
          12'h833: exp_out = 32'h00000168; // x = -15.6016, f(x) = 0.0000
          12'h834: exp_out = 32'h0000016B; // x = -15.5938, f(x) = 0.0000
          12'h835: exp_out = 32'h0000016E; // x = -15.5859, f(x) = 0.0000
          12'h836: exp_out = 32'h00000170; // x = -15.5781, f(x) = 0.0000
          12'h837: exp_out = 32'h00000173; // x = -15.5703, f(x) = 0.0000
          12'h838: exp_out = 32'h00000176; // x = -15.5625, f(x) = 0.0000
          12'h839: exp_out = 32'h00000179; // x = -15.5547, f(x) = 0.0000
          12'h83A: exp_out = 32'h0000017C; // x = -15.5469, f(x) = 0.0000
          12'h83B: exp_out = 32'h0000017F; // x = -15.5391, f(x) = 0.0000
          12'h83C: exp_out = 32'h00000182; // x = -15.5312, f(x) = 0.0000
          12'h83D: exp_out = 32'h00000185; // x = -15.5234, f(x) = 0.0000
          12'h83E: exp_out = 32'h00000188; // x = -15.5156, f(x) = 0.0000
          12'h83F: exp_out = 32'h0000018B; // x = -15.5078, f(x) = 0.0000
          12'h840: exp_out = 32'h0000018E; // x = -15.5000, f(x) = 0.0000
          12'h841: exp_out = 32'h00000192; // x = -15.4922, f(x) = 0.0000
          12'h842: exp_out = 32'h00000195; // x = -15.4844, f(x) = 0.0000
          12'h843: exp_out = 32'h00000198; // x = -15.4766, f(x) = 0.0000
          12'h844: exp_out = 32'h0000019B; // x = -15.4688, f(x) = 0.0000
          12'h845: exp_out = 32'h0000019E; // x = -15.4609, f(x) = 0.0000
          12'h846: exp_out = 32'h000001A2; // x = -15.4531, f(x) = 0.0000
          12'h847: exp_out = 32'h000001A5; // x = -15.4453, f(x) = 0.0000
          12'h848: exp_out = 32'h000001A8; // x = -15.4375, f(x) = 0.0000
          12'h849: exp_out = 32'h000001AB; // x = -15.4297, f(x) = 0.0000
          12'h84A: exp_out = 32'h000001AF; // x = -15.4219, f(x) = 0.0000
          12'h84B: exp_out = 32'h000001B2; // x = -15.4141, f(x) = 0.0000
          12'h84C: exp_out = 32'h000001B6; // x = -15.4062, f(x) = 0.0000
          12'h84D: exp_out = 32'h000001B9; // x = -15.3984, f(x) = 0.0000
          12'h84E: exp_out = 32'h000001BC; // x = -15.3906, f(x) = 0.0000
          12'h84F: exp_out = 32'h000001C0; // x = -15.3828, f(x) = 0.0000
          12'h850: exp_out = 32'h000001C3; // x = -15.3750, f(x) = 0.0000
          12'h851: exp_out = 32'h000001C7; // x = -15.3672, f(x) = 0.0000
          12'h852: exp_out = 32'h000001CB; // x = -15.3594, f(x) = 0.0000
          12'h853: exp_out = 32'h000001CE; // x = -15.3516, f(x) = 0.0000
          12'h854: exp_out = 32'h000001D2; // x = -15.3438, f(x) = 0.0000
          12'h855: exp_out = 32'h000001D5; // x = -15.3359, f(x) = 0.0000
          12'h856: exp_out = 32'h000001D9; // x = -15.3281, f(x) = 0.0000
          12'h857: exp_out = 32'h000001DD; // x = -15.3203, f(x) = 0.0000
          12'h858: exp_out = 32'h000001E1; // x = -15.3125, f(x) = 0.0000
          12'h859: exp_out = 32'h000001E4; // x = -15.3047, f(x) = 0.0000
          12'h85A: exp_out = 32'h000001E8; // x = -15.2969, f(x) = 0.0000
          12'h85B: exp_out = 32'h000001EC; // x = -15.2891, f(x) = 0.0000
          12'h85C: exp_out = 32'h000001F0; // x = -15.2812, f(x) = 0.0000
          12'h85D: exp_out = 32'h000001F4; // x = -15.2734, f(x) = 0.0000
          12'h85E: exp_out = 32'h000001F8; // x = -15.2656, f(x) = 0.0000
          12'h85F: exp_out = 32'h000001FC; // x = -15.2578, f(x) = 0.0000
          12'h860: exp_out = 32'h00000200; // x = -15.2500, f(x) = 0.0000
          12'h861: exp_out = 32'h00000204; // x = -15.2422, f(x) = 0.0000
          12'h862: exp_out = 32'h00000208; // x = -15.2344, f(x) = 0.0000
          12'h863: exp_out = 32'h0000020C; // x = -15.2266, f(x) = 0.0000
          12'h864: exp_out = 32'h00000210; // x = -15.2188, f(x) = 0.0000
          12'h865: exp_out = 32'h00000214; // x = -15.2109, f(x) = 0.0000
          12'h866: exp_out = 32'h00000218; // x = -15.2031, f(x) = 0.0000
          12'h867: exp_out = 32'h0000021C; // x = -15.1953, f(x) = 0.0000
          12'h868: exp_out = 32'h00000221; // x = -15.1875, f(x) = 0.0000
          12'h869: exp_out = 32'h00000225; // x = -15.1797, f(x) = 0.0000
          12'h86A: exp_out = 32'h00000229; // x = -15.1719, f(x) = 0.0000
          12'h86B: exp_out = 32'h0000022E; // x = -15.1641, f(x) = 0.0000
          12'h86C: exp_out = 32'h00000232; // x = -15.1562, f(x) = 0.0000
          12'h86D: exp_out = 32'h00000236; // x = -15.1484, f(x) = 0.0000
          12'h86E: exp_out = 32'h0000023B; // x = -15.1406, f(x) = 0.0000
          12'h86F: exp_out = 32'h0000023F; // x = -15.1328, f(x) = 0.0000
          12'h870: exp_out = 32'h00000244; // x = -15.1250, f(x) = 0.0000
          12'h871: exp_out = 32'h00000248; // x = -15.1172, f(x) = 0.0000
          12'h872: exp_out = 32'h0000024D; // x = -15.1094, f(x) = 0.0000
          12'h873: exp_out = 32'h00000251; // x = -15.1016, f(x) = 0.0000
          12'h874: exp_out = 32'h00000256; // x = -15.0938, f(x) = 0.0000
          12'h875: exp_out = 32'h0000025B; // x = -15.0859, f(x) = 0.0000
          12'h876: exp_out = 32'h00000260; // x = -15.0781, f(x) = 0.0000
          12'h877: exp_out = 32'h00000264; // x = -15.0703, f(x) = 0.0000
          12'h878: exp_out = 32'h00000269; // x = -15.0625, f(x) = 0.0000
          12'h879: exp_out = 32'h0000026E; // x = -15.0547, f(x) = 0.0000
          12'h87A: exp_out = 32'h00000273; // x = -15.0469, f(x) = 0.0000
          12'h87B: exp_out = 32'h00000278; // x = -15.0391, f(x) = 0.0000
          12'h87C: exp_out = 32'h0000027D; // x = -15.0312, f(x) = 0.0000
          12'h87D: exp_out = 32'h00000282; // x = -15.0234, f(x) = 0.0000
          12'h87E: exp_out = 32'h00000287; // x = -15.0156, f(x) = 0.0000
          12'h87F: exp_out = 32'h0000028C; // x = -15.0078, f(x) = 0.0000
          12'h880: exp_out = 32'h00000291; // x = -15.0000, f(x) = 0.0000
          12'h881: exp_out = 32'h00000296; // x = -14.9922, f(x) = 0.0000
          12'h882: exp_out = 32'h0000029B; // x = -14.9844, f(x) = 0.0000
          12'h883: exp_out = 32'h000002A0; // x = -14.9766, f(x) = 0.0000
          12'h884: exp_out = 32'h000002A6; // x = -14.9688, f(x) = 0.0000
          12'h885: exp_out = 32'h000002AB; // x = -14.9609, f(x) = 0.0000
          12'h886: exp_out = 32'h000002B0; // x = -14.9531, f(x) = 0.0000
          12'h887: exp_out = 32'h000002B6; // x = -14.9453, f(x) = 0.0000
          12'h888: exp_out = 32'h000002BB; // x = -14.9375, f(x) = 0.0000
          12'h889: exp_out = 32'h000002C1; // x = -14.9297, f(x) = 0.0000
          12'h88A: exp_out = 32'h000002C6; // x = -14.9219, f(x) = 0.0000
          12'h88B: exp_out = 32'h000002CC; // x = -14.9141, f(x) = 0.0000
          12'h88C: exp_out = 32'h000002D1; // x = -14.9062, f(x) = 0.0000
          12'h88D: exp_out = 32'h000002D7; // x = -14.8984, f(x) = 0.0000
          12'h88E: exp_out = 32'h000002DD; // x = -14.8906, f(x) = 0.0000
          12'h88F: exp_out = 32'h000002E3; // x = -14.8828, f(x) = 0.0000
          12'h890: exp_out = 32'h000002E8; // x = -14.8750, f(x) = 0.0000
          12'h891: exp_out = 32'h000002EE; // x = -14.8672, f(x) = 0.0000
          12'h892: exp_out = 32'h000002F4; // x = -14.8594, f(x) = 0.0000
          12'h893: exp_out = 32'h000002FA; // x = -14.8516, f(x) = 0.0000
          12'h894: exp_out = 32'h00000300; // x = -14.8438, f(x) = 0.0000
          12'h895: exp_out = 32'h00000306; // x = -14.8359, f(x) = 0.0000
          12'h896: exp_out = 32'h0000030C; // x = -14.8281, f(x) = 0.0000
          12'h897: exp_out = 32'h00000312; // x = -14.8203, f(x) = 0.0000
          12'h898: exp_out = 32'h00000318; // x = -14.8125, f(x) = 0.0000
          12'h899: exp_out = 32'h0000031F; // x = -14.8047, f(x) = 0.0000
          12'h89A: exp_out = 32'h00000325; // x = -14.7969, f(x) = 0.0000
          12'h89B: exp_out = 32'h0000032B; // x = -14.7891, f(x) = 0.0000
          12'h89C: exp_out = 32'h00000332; // x = -14.7812, f(x) = 0.0000
          12'h89D: exp_out = 32'h00000338; // x = -14.7734, f(x) = 0.0000
          12'h89E: exp_out = 32'h0000033E; // x = -14.7656, f(x) = 0.0000
          12'h89F: exp_out = 32'h00000345; // x = -14.7578, f(x) = 0.0000
          12'h8A0: exp_out = 32'h0000034C; // x = -14.7500, f(x) = 0.0000
          12'h8A1: exp_out = 32'h00000352; // x = -14.7422, f(x) = 0.0000
          12'h8A2: exp_out = 32'h00000359; // x = -14.7344, f(x) = 0.0000
          12'h8A3: exp_out = 32'h00000360; // x = -14.7266, f(x) = 0.0000
          12'h8A4: exp_out = 32'h00000366; // x = -14.7188, f(x) = 0.0000
          12'h8A5: exp_out = 32'h0000036D; // x = -14.7109, f(x) = 0.0000
          12'h8A6: exp_out = 32'h00000374; // x = -14.7031, f(x) = 0.0000
          12'h8A7: exp_out = 32'h0000037B; // x = -14.6953, f(x) = 0.0000
          12'h8A8: exp_out = 32'h00000382; // x = -14.6875, f(x) = 0.0000
          12'h8A9: exp_out = 32'h00000389; // x = -14.6797, f(x) = 0.0000
          12'h8AA: exp_out = 32'h00000390; // x = -14.6719, f(x) = 0.0000
          12'h8AB: exp_out = 32'h00000397; // x = -14.6641, f(x) = 0.0000
          12'h8AC: exp_out = 32'h0000039E; // x = -14.6562, f(x) = 0.0000
          12'h8AD: exp_out = 32'h000003A6; // x = -14.6484, f(x) = 0.0000
          12'h8AE: exp_out = 32'h000003AD; // x = -14.6406, f(x) = 0.0000
          12'h8AF: exp_out = 32'h000003B4; // x = -14.6328, f(x) = 0.0000
          12'h8B0: exp_out = 32'h000003BC; // x = -14.6250, f(x) = 0.0000
          12'h8B1: exp_out = 32'h000003C3; // x = -14.6172, f(x) = 0.0000
          12'h8B2: exp_out = 32'h000003CB; // x = -14.6094, f(x) = 0.0000
          12'h8B3: exp_out = 32'h000003D2; // x = -14.6016, f(x) = 0.0000
          12'h8B4: exp_out = 32'h000003DA; // x = -14.5938, f(x) = 0.0000
          12'h8B5: exp_out = 32'h000003E2; // x = -14.5859, f(x) = 0.0000
          12'h8B6: exp_out = 32'h000003EA; // x = -14.5781, f(x) = 0.0000
          12'h8B7: exp_out = 32'h000003F2; // x = -14.5703, f(x) = 0.0000
          12'h8B8: exp_out = 32'h000003F9; // x = -14.5625, f(x) = 0.0000
          12'h8B9: exp_out = 32'h00000401; // x = -14.5547, f(x) = 0.0000
          12'h8BA: exp_out = 32'h00000409; // x = -14.5469, f(x) = 0.0000
          12'h8BB: exp_out = 32'h00000412; // x = -14.5391, f(x) = 0.0000
          12'h8BC: exp_out = 32'h0000041A; // x = -14.5312, f(x) = 0.0000
          12'h8BD: exp_out = 32'h00000422; // x = -14.5234, f(x) = 0.0000
          12'h8BE: exp_out = 32'h0000042A; // x = -14.5156, f(x) = 0.0000
          12'h8BF: exp_out = 32'h00000433; // x = -14.5078, f(x) = 0.0000
          12'h8C0: exp_out = 32'h0000043B; // x = -14.5000, f(x) = 0.0000
          12'h8C1: exp_out = 32'h00000444; // x = -14.4922, f(x) = 0.0000
          12'h8C2: exp_out = 32'h0000044C; // x = -14.4844, f(x) = 0.0000
          12'h8C3: exp_out = 32'h00000455; // x = -14.4766, f(x) = 0.0000
          12'h8C4: exp_out = 32'h0000045D; // x = -14.4688, f(x) = 0.0000
          12'h8C5: exp_out = 32'h00000466; // x = -14.4609, f(x) = 0.0000
          12'h8C6: exp_out = 32'h0000046F; // x = -14.4531, f(x) = 0.0000
          12'h8C7: exp_out = 32'h00000478; // x = -14.4453, f(x) = 0.0000
          12'h8C8: exp_out = 32'h00000481; // x = -14.4375, f(x) = 0.0000
          12'h8C9: exp_out = 32'h0000048A; // x = -14.4297, f(x) = 0.0000
          12'h8CA: exp_out = 32'h00000493; // x = -14.4219, f(x) = 0.0000
          12'h8CB: exp_out = 32'h0000049C; // x = -14.4141, f(x) = 0.0000
          12'h8CC: exp_out = 32'h000004A6; // x = -14.4062, f(x) = 0.0000
          12'h8CD: exp_out = 32'h000004AF; // x = -14.3984, f(x) = 0.0000
          12'h8CE: exp_out = 32'h000004B8; // x = -14.3906, f(x) = 0.0000
          12'h8CF: exp_out = 32'h000004C2; // x = -14.3828, f(x) = 0.0000
          12'h8D0: exp_out = 32'h000004CB; // x = -14.3750, f(x) = 0.0000
          12'h8D1: exp_out = 32'h000004D5; // x = -14.3672, f(x) = 0.0000
          12'h8D2: exp_out = 32'h000004DF; // x = -14.3594, f(x) = 0.0000
          12'h8D3: exp_out = 32'h000004E8; // x = -14.3516, f(x) = 0.0000
          12'h8D4: exp_out = 32'h000004F2; // x = -14.3438, f(x) = 0.0000
          12'h8D5: exp_out = 32'h000004FC; // x = -14.3359, f(x) = 0.0000
          12'h8D6: exp_out = 32'h00000506; // x = -14.3281, f(x) = 0.0000
          12'h8D7: exp_out = 32'h00000510; // x = -14.3203, f(x) = 0.0000
          12'h8D8: exp_out = 32'h0000051A; // x = -14.3125, f(x) = 0.0000
          12'h8D9: exp_out = 32'h00000525; // x = -14.3047, f(x) = 0.0000
          12'h8DA: exp_out = 32'h0000052F; // x = -14.2969, f(x) = 0.0000
          12'h8DB: exp_out = 32'h00000539; // x = -14.2891, f(x) = 0.0000
          12'h8DC: exp_out = 32'h00000544; // x = -14.2812, f(x) = 0.0000
          12'h8DD: exp_out = 32'h0000054E; // x = -14.2734, f(x) = 0.0000
          12'h8DE: exp_out = 32'h00000559; // x = -14.2656, f(x) = 0.0000
          12'h8DF: exp_out = 32'h00000564; // x = -14.2578, f(x) = 0.0000
          12'h8E0: exp_out = 32'h0000056F; // x = -14.2500, f(x) = 0.0000
          12'h8E1: exp_out = 32'h0000057A; // x = -14.2422, f(x) = 0.0000
          12'h8E2: exp_out = 32'h00000585; // x = -14.2344, f(x) = 0.0000
          12'h8E3: exp_out = 32'h00000590; // x = -14.2266, f(x) = 0.0000
          12'h8E4: exp_out = 32'h0000059B; // x = -14.2188, f(x) = 0.0000
          12'h8E5: exp_out = 32'h000005A6; // x = -14.2109, f(x) = 0.0000
          12'h8E6: exp_out = 32'h000005B1; // x = -14.2031, f(x) = 0.0000
          12'h8E7: exp_out = 32'h000005BD; // x = -14.1953, f(x) = 0.0000
          12'h8E8: exp_out = 32'h000005C8; // x = -14.1875, f(x) = 0.0000
          12'h8E9: exp_out = 32'h000005D4; // x = -14.1797, f(x) = 0.0000
          12'h8EA: exp_out = 32'h000005E0; // x = -14.1719, f(x) = 0.0000
          12'h8EB: exp_out = 32'h000005EB; // x = -14.1641, f(x) = 0.0000
          12'h8EC: exp_out = 32'h000005F7; // x = -14.1562, f(x) = 0.0000
          12'h8ED: exp_out = 32'h00000603; // x = -14.1484, f(x) = 0.0000
          12'h8EE: exp_out = 32'h0000060F; // x = -14.1406, f(x) = 0.0000
          12'h8EF: exp_out = 32'h0000061C; // x = -14.1328, f(x) = 0.0000
          12'h8F0: exp_out = 32'h00000628; // x = -14.1250, f(x) = 0.0000
          12'h8F1: exp_out = 32'h00000634; // x = -14.1172, f(x) = 0.0000
          12'h8F2: exp_out = 32'h00000641; // x = -14.1094, f(x) = 0.0000
          12'h8F3: exp_out = 32'h0000064D; // x = -14.1016, f(x) = 0.0000
          12'h8F4: exp_out = 32'h0000065A; // x = -14.0938, f(x) = 0.0000
          12'h8F5: exp_out = 32'h00000667; // x = -14.0859, f(x) = 0.0000
          12'h8F6: exp_out = 32'h00000673; // x = -14.0781, f(x) = 0.0000
          12'h8F7: exp_out = 32'h00000680; // x = -14.0703, f(x) = 0.0000
          12'h8F8: exp_out = 32'h0000068E; // x = -14.0625, f(x) = 0.0000
          12'h8F9: exp_out = 32'h0000069B; // x = -14.0547, f(x) = 0.0000
          12'h8FA: exp_out = 32'h000006A8; // x = -14.0469, f(x) = 0.0000
          12'h8FB: exp_out = 32'h000006B5; // x = -14.0391, f(x) = 0.0000
          12'h8FC: exp_out = 32'h000006C3; // x = -14.0312, f(x) = 0.0000
          12'h8FD: exp_out = 32'h000006D0; // x = -14.0234, f(x) = 0.0000
          12'h8FE: exp_out = 32'h000006DE; // x = -14.0156, f(x) = 0.0000
          12'h8FF: exp_out = 32'h000006EC; // x = -14.0078, f(x) = 0.0000
          12'h900: exp_out = 32'h000006FA; // x = -14.0000, f(x) = 0.0000
          12'h901: exp_out = 32'h00000708; // x = -13.9922, f(x) = 0.0000
          12'h902: exp_out = 32'h00000716; // x = -13.9844, f(x) = 0.0000
          12'h903: exp_out = 32'h00000724; // x = -13.9766, f(x) = 0.0000
          12'h904: exp_out = 32'h00000732; // x = -13.9688, f(x) = 0.0000
          12'h905: exp_out = 32'h00000741; // x = -13.9609, f(x) = 0.0000
          12'h906: exp_out = 32'h0000074F; // x = -13.9531, f(x) = 0.0000
          12'h907: exp_out = 32'h0000075E; // x = -13.9453, f(x) = 0.0000
          12'h908: exp_out = 32'h0000076D; // x = -13.9375, f(x) = 0.0000
          12'h909: exp_out = 32'h0000077C; // x = -13.9297, f(x) = 0.0000
          12'h90A: exp_out = 32'h0000078B; // x = -13.9219, f(x) = 0.0000
          12'h90B: exp_out = 32'h0000079A; // x = -13.9141, f(x) = 0.0000
          12'h90C: exp_out = 32'h000007A9; // x = -13.9062, f(x) = 0.0000
          12'h90D: exp_out = 32'h000007B9; // x = -13.8984, f(x) = 0.0000
          12'h90E: exp_out = 32'h000007C8; // x = -13.8906, f(x) = 0.0000
          12'h90F: exp_out = 32'h000007D8; // x = -13.8828, f(x) = 0.0000
          12'h910: exp_out = 32'h000007E7; // x = -13.8750, f(x) = 0.0000
          12'h911: exp_out = 32'h000007F7; // x = -13.8672, f(x) = 0.0000
          12'h912: exp_out = 32'h00000807; // x = -13.8594, f(x) = 0.0000
          12'h913: exp_out = 32'h00000817; // x = -13.8516, f(x) = 0.0000
          12'h914: exp_out = 32'h00000828; // x = -13.8438, f(x) = 0.0000
          12'h915: exp_out = 32'h00000838; // x = -13.8359, f(x) = 0.0000
          12'h916: exp_out = 32'h00000849; // x = -13.8281, f(x) = 0.0000
          12'h917: exp_out = 32'h00000859; // x = -13.8203, f(x) = 0.0000
          12'h918: exp_out = 32'h0000086A; // x = -13.8125, f(x) = 0.0000
          12'h919: exp_out = 32'h0000087B; // x = -13.8047, f(x) = 0.0000
          12'h91A: exp_out = 32'h0000088C; // x = -13.7969, f(x) = 0.0000
          12'h91B: exp_out = 32'h0000089D; // x = -13.7891, f(x) = 0.0000
          12'h91C: exp_out = 32'h000008AE; // x = -13.7812, f(x) = 0.0000
          12'h91D: exp_out = 32'h000008C0; // x = -13.7734, f(x) = 0.0000
          12'h91E: exp_out = 32'h000008D1; // x = -13.7656, f(x) = 0.0000
          12'h91F: exp_out = 32'h000008E3; // x = -13.7578, f(x) = 0.0000
          12'h920: exp_out = 32'h000008F5; // x = -13.7500, f(x) = 0.0000
          12'h921: exp_out = 32'h00000907; // x = -13.7422, f(x) = 0.0000
          12'h922: exp_out = 32'h00000919; // x = -13.7344, f(x) = 0.0000
          12'h923: exp_out = 32'h0000092B; // x = -13.7266, f(x) = 0.0000
          12'h924: exp_out = 32'h0000093E; // x = -13.7188, f(x) = 0.0000
          12'h925: exp_out = 32'h00000950; // x = -13.7109, f(x) = 0.0000
          12'h926: exp_out = 32'h00000963; // x = -13.7031, f(x) = 0.0000
          12'h927: exp_out = 32'h00000976; // x = -13.6953, f(x) = 0.0000
          12'h928: exp_out = 32'h00000989; // x = -13.6875, f(x) = 0.0000
          12'h929: exp_out = 32'h0000099C; // x = -13.6797, f(x) = 0.0000
          12'h92A: exp_out = 32'h000009AF; // x = -13.6719, f(x) = 0.0000
          12'h92B: exp_out = 32'h000009C3; // x = -13.6641, f(x) = 0.0000
          12'h92C: exp_out = 32'h000009D6; // x = -13.6562, f(x) = 0.0000
          12'h92D: exp_out = 32'h000009EA; // x = -13.6484, f(x) = 0.0000
          12'h92E: exp_out = 32'h000009FE; // x = -13.6406, f(x) = 0.0000
          12'h92F: exp_out = 32'h00000A12; // x = -13.6328, f(x) = 0.0000
          12'h930: exp_out = 32'h00000A26; // x = -13.6250, f(x) = 0.0000
          12'h931: exp_out = 32'h00000A3B; // x = -13.6172, f(x) = 0.0000
          12'h932: exp_out = 32'h00000A4F; // x = -13.6094, f(x) = 0.0000
          12'h933: exp_out = 32'h00000A64; // x = -13.6016, f(x) = 0.0000
          12'h934: exp_out = 32'h00000A79; // x = -13.5938, f(x) = 0.0000
          12'h935: exp_out = 32'h00000A8E; // x = -13.5859, f(x) = 0.0000
          12'h936: exp_out = 32'h00000AA3; // x = -13.5781, f(x) = 0.0000
          12'h937: exp_out = 32'h00000AB8; // x = -13.5703, f(x) = 0.0000
          12'h938: exp_out = 32'h00000ACE; // x = -13.5625, f(x) = 0.0000
          12'h939: exp_out = 32'h00000AE3; // x = -13.5547, f(x) = 0.0000
          12'h93A: exp_out = 32'h00000AF9; // x = -13.5469, f(x) = 0.0000
          12'h93B: exp_out = 32'h00000B0F; // x = -13.5391, f(x) = 0.0000
          12'h93C: exp_out = 32'h00000B26; // x = -13.5312, f(x) = 0.0000
          12'h93D: exp_out = 32'h00000B3C; // x = -13.5234, f(x) = 0.0000
          12'h93E: exp_out = 32'h00000B52; // x = -13.5156, f(x) = 0.0000
          12'h93F: exp_out = 32'h00000B69; // x = -13.5078, f(x) = 0.0000
          12'h940: exp_out = 32'h00000B80; // x = -13.5000, f(x) = 0.0000
          12'h941: exp_out = 32'h00000B97; // x = -13.4922, f(x) = 0.0000
          12'h942: exp_out = 32'h00000BAE; // x = -13.4844, f(x) = 0.0000
          12'h943: exp_out = 32'h00000BC6; // x = -13.4766, f(x) = 0.0000
          12'h944: exp_out = 32'h00000BDE; // x = -13.4688, f(x) = 0.0000
          12'h945: exp_out = 32'h00000BF5; // x = -13.4609, f(x) = 0.0000
          12'h946: exp_out = 32'h00000C0D; // x = -13.4531, f(x) = 0.0000
          12'h947: exp_out = 32'h00000C26; // x = -13.4453, f(x) = 0.0000
          12'h948: exp_out = 32'h00000C3E; // x = -13.4375, f(x) = 0.0000
          12'h949: exp_out = 32'h00000C57; // x = -13.4297, f(x) = 0.0000
          12'h94A: exp_out = 32'h00000C6F; // x = -13.4219, f(x) = 0.0000
          12'h94B: exp_out = 32'h00000C88; // x = -13.4141, f(x) = 0.0000
          12'h94C: exp_out = 32'h00000CA1; // x = -13.4062, f(x) = 0.0000
          12'h94D: exp_out = 32'h00000CBB; // x = -13.3984, f(x) = 0.0000
          12'h94E: exp_out = 32'h00000CD4; // x = -13.3906, f(x) = 0.0000
          12'h94F: exp_out = 32'h00000CEE; // x = -13.3828, f(x) = 0.0000
          12'h950: exp_out = 32'h00000D08; // x = -13.3750, f(x) = 0.0000
          12'h951: exp_out = 32'h00000D22; // x = -13.3672, f(x) = 0.0000
          12'h952: exp_out = 32'h00000D3D; // x = -13.3594, f(x) = 0.0000
          12'h953: exp_out = 32'h00000D57; // x = -13.3516, f(x) = 0.0000
          12'h954: exp_out = 32'h00000D72; // x = -13.3438, f(x) = 0.0000
          12'h955: exp_out = 32'h00000D8D; // x = -13.3359, f(x) = 0.0000
          12'h956: exp_out = 32'h00000DA8; // x = -13.3281, f(x) = 0.0000
          12'h957: exp_out = 32'h00000DC4; // x = -13.3203, f(x) = 0.0000
          12'h958: exp_out = 32'h00000DDF; // x = -13.3125, f(x) = 0.0000
          12'h959: exp_out = 32'h00000DFB; // x = -13.3047, f(x) = 0.0000
          12'h95A: exp_out = 32'h00000E17; // x = -13.2969, f(x) = 0.0000
          12'h95B: exp_out = 32'h00000E33; // x = -13.2891, f(x) = 0.0000
          12'h95C: exp_out = 32'h00000E50; // x = -13.2812, f(x) = 0.0000
          12'h95D: exp_out = 32'h00000E6D; // x = -13.2734, f(x) = 0.0000
          12'h95E: exp_out = 32'h00000E8A; // x = -13.2656, f(x) = 0.0000
          12'h95F: exp_out = 32'h00000EA7; // x = -13.2578, f(x) = 0.0000
          12'h960: exp_out = 32'h00000EC4; // x = -13.2500, f(x) = 0.0000
          12'h961: exp_out = 32'h00000EE2; // x = -13.2422, f(x) = 0.0000
          12'h962: exp_out = 32'h00000F00; // x = -13.2344, f(x) = 0.0000
          12'h963: exp_out = 32'h00000F1E; // x = -13.2266, f(x) = 0.0000
          12'h964: exp_out = 32'h00000F3C; // x = -13.2188, f(x) = 0.0000
          12'h965: exp_out = 32'h00000F5B; // x = -13.2109, f(x) = 0.0000
          12'h966: exp_out = 32'h00000F7A; // x = -13.2031, f(x) = 0.0000
          12'h967: exp_out = 32'h00000F99; // x = -13.1953, f(x) = 0.0000
          12'h968: exp_out = 32'h00000FB8; // x = -13.1875, f(x) = 0.0000
          12'h969: exp_out = 32'h00000FD8; // x = -13.1797, f(x) = 0.0000
          12'h96A: exp_out = 32'h00000FF7; // x = -13.1719, f(x) = 0.0000
          12'h96B: exp_out = 32'h00001018; // x = -13.1641, f(x) = 0.0000
          12'h96C: exp_out = 32'h00001038; // x = -13.1562, f(x) = 0.0000
          12'h96D: exp_out = 32'h00001058; // x = -13.1484, f(x) = 0.0000
          12'h96E: exp_out = 32'h00001079; // x = -13.1406, f(x) = 0.0000
          12'h96F: exp_out = 32'h0000109A; // x = -13.1328, f(x) = 0.0000
          12'h970: exp_out = 32'h000010BC; // x = -13.1250, f(x) = 0.0000
          12'h971: exp_out = 32'h000010DD; // x = -13.1172, f(x) = 0.0000
          12'h972: exp_out = 32'h000010FF; // x = -13.1094, f(x) = 0.0000
          12'h973: exp_out = 32'h00001121; // x = -13.1016, f(x) = 0.0000
          12'h974: exp_out = 32'h00001144; // x = -13.0938, f(x) = 0.0000
          12'h975: exp_out = 32'h00001166; // x = -13.0859, f(x) = 0.0000
          12'h976: exp_out = 32'h00001189; // x = -13.0781, f(x) = 0.0000
          12'h977: exp_out = 32'h000011AC; // x = -13.0703, f(x) = 0.0000
          12'h978: exp_out = 32'h000011D0; // x = -13.0625, f(x) = 0.0000
          12'h979: exp_out = 32'h000011F4; // x = -13.0547, f(x) = 0.0000
          12'h97A: exp_out = 32'h00001218; // x = -13.0469, f(x) = 0.0000
          12'h97B: exp_out = 32'h0000123C; // x = -13.0391, f(x) = 0.0000
          12'h97C: exp_out = 32'h00001261; // x = -13.0312, f(x) = 0.0000
          12'h97D: exp_out = 32'h00001286; // x = -13.0234, f(x) = 0.0000
          12'h97E: exp_out = 32'h000012AB; // x = -13.0156, f(x) = 0.0000
          12'h97F: exp_out = 32'h000012D0; // x = -13.0078, f(x) = 0.0000
          12'h980: exp_out = 32'h000012F6; // x = -13.0000, f(x) = 0.0000
          12'h981: exp_out = 32'h0000131C; // x = -12.9922, f(x) = 0.0000
          12'h982: exp_out = 32'h00001342; // x = -12.9844, f(x) = 0.0000
          12'h983: exp_out = 32'h00001369; // x = -12.9766, f(x) = 0.0000
          12'h984: exp_out = 32'h00001390; // x = -12.9688, f(x) = 0.0000
          12'h985: exp_out = 32'h000013B7; // x = -12.9609, f(x) = 0.0000
          12'h986: exp_out = 32'h000013DF; // x = -12.9531, f(x) = 0.0000
          12'h987: exp_out = 32'h00001407; // x = -12.9453, f(x) = 0.0000
          12'h988: exp_out = 32'h0000142F; // x = -12.9375, f(x) = 0.0000
          12'h989: exp_out = 32'h00001458; // x = -12.9297, f(x) = 0.0000
          12'h98A: exp_out = 32'h00001480; // x = -12.9219, f(x) = 0.0000
          12'h98B: exp_out = 32'h000014AA; // x = -12.9141, f(x) = 0.0000
          12'h98C: exp_out = 32'h000014D3; // x = -12.9062, f(x) = 0.0000
          12'h98D: exp_out = 32'h000014FD; // x = -12.8984, f(x) = 0.0000
          12'h98E: exp_out = 32'h00001527; // x = -12.8906, f(x) = 0.0000
          12'h98F: exp_out = 32'h00001552; // x = -12.8828, f(x) = 0.0000
          12'h990: exp_out = 32'h0000157C; // x = -12.8750, f(x) = 0.0000
          12'h991: exp_out = 32'h000015A7; // x = -12.8672, f(x) = 0.0000
          12'h992: exp_out = 32'h000015D3; // x = -12.8594, f(x) = 0.0000
          12'h993: exp_out = 32'h000015FF; // x = -12.8516, f(x) = 0.0000
          12'h994: exp_out = 32'h0000162B; // x = -12.8438, f(x) = 0.0000
          12'h995: exp_out = 32'h00001657; // x = -12.8359, f(x) = 0.0000
          12'h996: exp_out = 32'h00001684; // x = -12.8281, f(x) = 0.0000
          12'h997: exp_out = 32'h000016B2; // x = -12.8203, f(x) = 0.0000
          12'h998: exp_out = 32'h000016DF; // x = -12.8125, f(x) = 0.0000
          12'h999: exp_out = 32'h0000170D; // x = -12.8047, f(x) = 0.0000
          12'h99A: exp_out = 32'h0000173B; // x = -12.7969, f(x) = 0.0000
          12'h99B: exp_out = 32'h0000176A; // x = -12.7891, f(x) = 0.0000
          12'h99C: exp_out = 32'h00001799; // x = -12.7812, f(x) = 0.0000
          12'h99D: exp_out = 32'h000017C8; // x = -12.7734, f(x) = 0.0000
          12'h99E: exp_out = 32'h000017F8; // x = -12.7656, f(x) = 0.0000
          12'h99F: exp_out = 32'h00001828; // x = -12.7578, f(x) = 0.0000
          12'h9A0: exp_out = 32'h00001859; // x = -12.7500, f(x) = 0.0000
          12'h9A1: exp_out = 32'h0000188A; // x = -12.7422, f(x) = 0.0000
          12'h9A2: exp_out = 32'h000018BB; // x = -12.7344, f(x) = 0.0000
          12'h9A3: exp_out = 32'h000018EC; // x = -12.7266, f(x) = 0.0000
          12'h9A4: exp_out = 32'h0000191F; // x = -12.7188, f(x) = 0.0000
          12'h9A5: exp_out = 32'h00001951; // x = -12.7109, f(x) = 0.0000
          12'h9A6: exp_out = 32'h00001984; // x = -12.7031, f(x) = 0.0000
          12'h9A7: exp_out = 32'h000019B7; // x = -12.6953, f(x) = 0.0000
          12'h9A8: exp_out = 32'h000019EB; // x = -12.6875, f(x) = 0.0000
          12'h9A9: exp_out = 32'h00001A1F; // x = -12.6797, f(x) = 0.0000
          12'h9AA: exp_out = 32'h00001A53; // x = -12.6719, f(x) = 0.0000
          12'h9AB: exp_out = 32'h00001A88; // x = -12.6641, f(x) = 0.0000
          12'h9AC: exp_out = 32'h00001ABD; // x = -12.6562, f(x) = 0.0000
          12'h9AD: exp_out = 32'h00001AF3; // x = -12.6484, f(x) = 0.0000
          12'h9AE: exp_out = 32'h00001B29; // x = -12.6406, f(x) = 0.0000
          12'h9AF: exp_out = 32'h00001B60; // x = -12.6328, f(x) = 0.0000
          12'h9B0: exp_out = 32'h00001B97; // x = -12.6250, f(x) = 0.0000
          12'h9B1: exp_out = 32'h00001BCE; // x = -12.6172, f(x) = 0.0000
          12'h9B2: exp_out = 32'h00001C06; // x = -12.6094, f(x) = 0.0000
          12'h9B3: exp_out = 32'h00001C3E; // x = -12.6016, f(x) = 0.0000
          12'h9B4: exp_out = 32'h00001C77; // x = -12.5938, f(x) = 0.0000
          12'h9B5: exp_out = 32'h00001CB0; // x = -12.5859, f(x) = 0.0000
          12'h9B6: exp_out = 32'h00001CE9; // x = -12.5781, f(x) = 0.0000
          12'h9B7: exp_out = 32'h00001D24; // x = -12.5703, f(x) = 0.0000
          12'h9B8: exp_out = 32'h00001D5E; // x = -12.5625, f(x) = 0.0000
          12'h9B9: exp_out = 32'h00001D99; // x = -12.5547, f(x) = 0.0000
          12'h9BA: exp_out = 32'h00001DD4; // x = -12.5469, f(x) = 0.0000
          12'h9BB: exp_out = 32'h00001E10; // x = -12.5391, f(x) = 0.0000
          12'h9BC: exp_out = 32'h00001E4D; // x = -12.5312, f(x) = 0.0000
          12'h9BD: exp_out = 32'h00001E8A; // x = -12.5234, f(x) = 0.0000
          12'h9BE: exp_out = 32'h00001EC7; // x = -12.5156, f(x) = 0.0000
          12'h9BF: exp_out = 32'h00001F05; // x = -12.5078, f(x) = 0.0000
          12'h9C0: exp_out = 32'h00001F43; // x = -12.5000, f(x) = 0.0000
          12'h9C1: exp_out = 32'h00001F82; // x = -12.4922, f(x) = 0.0000
          12'h9C2: exp_out = 32'h00001FC1; // x = -12.4844, f(x) = 0.0000
          12'h9C3: exp_out = 32'h00002001; // x = -12.4766, f(x) = 0.0000
          12'h9C4: exp_out = 32'h00002041; // x = -12.4688, f(x) = 0.0000
          12'h9C5: exp_out = 32'h00002082; // x = -12.4609, f(x) = 0.0000
          12'h9C6: exp_out = 32'h000020C3; // x = -12.4531, f(x) = 0.0000
          12'h9C7: exp_out = 32'h00002105; // x = -12.4453, f(x) = 0.0000
          12'h9C8: exp_out = 32'h00002147; // x = -12.4375, f(x) = 0.0000
          12'h9C9: exp_out = 32'h0000218A; // x = -12.4297, f(x) = 0.0000
          12'h9CA: exp_out = 32'h000021CD; // x = -12.4219, f(x) = 0.0000
          12'h9CB: exp_out = 32'h00002211; // x = -12.4141, f(x) = 0.0000
          12'h9CC: exp_out = 32'h00002255; // x = -12.4062, f(x) = 0.0000
          12'h9CD: exp_out = 32'h0000229A; // x = -12.3984, f(x) = 0.0000
          12'h9CE: exp_out = 32'h000022E0; // x = -12.3906, f(x) = 0.0000
          12'h9CF: exp_out = 32'h00002326; // x = -12.3828, f(x) = 0.0000
          12'h9D0: exp_out = 32'h0000236D; // x = -12.3750, f(x) = 0.0000
          12'h9D1: exp_out = 32'h000023B4; // x = -12.3672, f(x) = 0.0000
          12'h9D2: exp_out = 32'h000023FB; // x = -12.3594, f(x) = 0.0000
          12'h9D3: exp_out = 32'h00002444; // x = -12.3516, f(x) = 0.0000
          12'h9D4: exp_out = 32'h0000248C; // x = -12.3438, f(x) = 0.0000
          12'h9D5: exp_out = 32'h000024D6; // x = -12.3359, f(x) = 0.0000
          12'h9D6: exp_out = 32'h00002520; // x = -12.3281, f(x) = 0.0000
          12'h9D7: exp_out = 32'h0000256A; // x = -12.3203, f(x) = 0.0000
          12'h9D8: exp_out = 32'h000025B5; // x = -12.3125, f(x) = 0.0000
          12'h9D9: exp_out = 32'h00002601; // x = -12.3047, f(x) = 0.0000
          12'h9DA: exp_out = 32'h0000264D; // x = -12.2969, f(x) = 0.0000
          12'h9DB: exp_out = 32'h0000269A; // x = -12.2891, f(x) = 0.0000
          12'h9DC: exp_out = 32'h000026E8; // x = -12.2812, f(x) = 0.0000
          12'h9DD: exp_out = 32'h00002736; // x = -12.2734, f(x) = 0.0000
          12'h9DE: exp_out = 32'h00002785; // x = -12.2656, f(x) = 0.0000
          12'h9DF: exp_out = 32'h000027D4; // x = -12.2578, f(x) = 0.0000
          12'h9E0: exp_out = 32'h00002824; // x = -12.2500, f(x) = 0.0000
          12'h9E1: exp_out = 32'h00002875; // x = -12.2422, f(x) = 0.0000
          12'h9E2: exp_out = 32'h000028C6; // x = -12.2344, f(x) = 0.0000
          12'h9E3: exp_out = 32'h00002918; // x = -12.2266, f(x) = 0.0000
          12'h9E4: exp_out = 32'h0000296A; // x = -12.2188, f(x) = 0.0000
          12'h9E5: exp_out = 32'h000029BD; // x = -12.2109, f(x) = 0.0000
          12'h9E6: exp_out = 32'h00002A11; // x = -12.2031, f(x) = 0.0000
          12'h9E7: exp_out = 32'h00002A66; // x = -12.1953, f(x) = 0.0000
          12'h9E8: exp_out = 32'h00002ABB; // x = -12.1875, f(x) = 0.0000
          12'h9E9: exp_out = 32'h00002B10; // x = -12.1797, f(x) = 0.0000
          12'h9EA: exp_out = 32'h00002B67; // x = -12.1719, f(x) = 0.0000
          12'h9EB: exp_out = 32'h00002BBE; // x = -12.1641, f(x) = 0.0000
          12'h9EC: exp_out = 32'h00002C16; // x = -12.1562, f(x) = 0.0000
          12'h9ED: exp_out = 32'h00002C6E; // x = -12.1484, f(x) = 0.0000
          12'h9EE: exp_out = 32'h00002CC8; // x = -12.1406, f(x) = 0.0000
          12'h9EF: exp_out = 32'h00002D22; // x = -12.1328, f(x) = 0.0000
          12'h9F0: exp_out = 32'h00002D7C; // x = -12.1250, f(x) = 0.0000
          12'h9F1: exp_out = 32'h00002DD8; // x = -12.1172, f(x) = 0.0000
          12'h9F2: exp_out = 32'h00002E34; // x = -12.1094, f(x) = 0.0000
          12'h9F3: exp_out = 32'h00002E90; // x = -12.1016, f(x) = 0.0000
          12'h9F4: exp_out = 32'h00002EEE; // x = -12.0938, f(x) = 0.0000
          12'h9F5: exp_out = 32'h00002F4C; // x = -12.0859, f(x) = 0.0000
          12'h9F6: exp_out = 32'h00002FAB; // x = -12.0781, f(x) = 0.0000
          12'h9F7: exp_out = 32'h0000300B; // x = -12.0703, f(x) = 0.0000
          12'h9F8: exp_out = 32'h0000306B; // x = -12.0625, f(x) = 0.0000
          12'h9F9: exp_out = 32'h000030CC; // x = -12.0547, f(x) = 0.0000
          12'h9FA: exp_out = 32'h0000312E; // x = -12.0469, f(x) = 0.0000
          12'h9FB: exp_out = 32'h00003191; // x = -12.0391, f(x) = 0.0000
          12'h9FC: exp_out = 32'h000031F5; // x = -12.0312, f(x) = 0.0000
          12'h9FD: exp_out = 32'h00003259; // x = -12.0234, f(x) = 0.0000
          12'h9FE: exp_out = 32'h000032BE; // x = -12.0156, f(x) = 0.0000
          12'h9FF: exp_out = 32'h00003324; // x = -12.0078, f(x) = 0.0000
          12'hA00: exp_out = 32'h0000338B; // x = -12.0000, f(x) = 0.0000
          12'hA01: exp_out = 32'h000033F2; // x = -11.9922, f(x) = 0.0000
          12'hA02: exp_out = 32'h0000345A; // x = -11.9844, f(x) = 0.0000
          12'hA03: exp_out = 32'h000034C3; // x = -11.9766, f(x) = 0.0000
          12'hA04: exp_out = 32'h0000352D; // x = -11.9688, f(x) = 0.0000
          12'hA05: exp_out = 32'h00003598; // x = -11.9609, f(x) = 0.0000
          12'hA06: exp_out = 32'h00003604; // x = -11.9531, f(x) = 0.0000
          12'hA07: exp_out = 32'h00003670; // x = -11.9453, f(x) = 0.0000
          12'hA08: exp_out = 32'h000036DE; // x = -11.9375, f(x) = 0.0000
          12'hA09: exp_out = 32'h0000374C; // x = -11.9297, f(x) = 0.0000
          12'hA0A: exp_out = 32'h000037BB; // x = -11.9219, f(x) = 0.0000
          12'hA0B: exp_out = 32'h0000382B; // x = -11.9141, f(x) = 0.0000
          12'hA0C: exp_out = 32'h0000389B; // x = -11.9062, f(x) = 0.0000
          12'hA0D: exp_out = 32'h0000390D; // x = -11.8984, f(x) = 0.0000
          12'hA0E: exp_out = 32'h00003980; // x = -11.8906, f(x) = 0.0000
          12'hA0F: exp_out = 32'h000039F3; // x = -11.8828, f(x) = 0.0000
          12'hA10: exp_out = 32'h00003A67; // x = -11.8750, f(x) = 0.0000
          12'hA11: exp_out = 32'h00003ADD; // x = -11.8672, f(x) = 0.0000
          12'hA12: exp_out = 32'h00003B53; // x = -11.8594, f(x) = 0.0000
          12'hA13: exp_out = 32'h00003BCA; // x = -11.8516, f(x) = 0.0000
          12'hA14: exp_out = 32'h00003C42; // x = -11.8438, f(x) = 0.0000
          12'hA15: exp_out = 32'h00003CBB; // x = -11.8359, f(x) = 0.0000
          12'hA16: exp_out = 32'h00003D35; // x = -11.8281, f(x) = 0.0000
          12'hA17: exp_out = 32'h00003DB0; // x = -11.8203, f(x) = 0.0000
          12'hA18: exp_out = 32'h00003E2C; // x = -11.8125, f(x) = 0.0000
          12'hA19: exp_out = 32'h00003EA9; // x = -11.8047, f(x) = 0.0000
          12'hA1A: exp_out = 32'h00003F26; // x = -11.7969, f(x) = 0.0000
          12'hA1B: exp_out = 32'h00003FA5; // x = -11.7891, f(x) = 0.0000
          12'hA1C: exp_out = 32'h00004025; // x = -11.7812, f(x) = 0.0000
          12'hA1D: exp_out = 32'h000040A6; // x = -11.7734, f(x) = 0.0000
          12'hA1E: exp_out = 32'h00004128; // x = -11.7656, f(x) = 0.0000
          12'hA1F: exp_out = 32'h000041AA; // x = -11.7578, f(x) = 0.0000
          12'hA20: exp_out = 32'h0000422E; // x = -11.7500, f(x) = 0.0000
          12'hA21: exp_out = 32'h000042B3; // x = -11.7422, f(x) = 0.0000
          12'hA22: exp_out = 32'h00004339; // x = -11.7344, f(x) = 0.0000
          12'hA23: exp_out = 32'h000043C0; // x = -11.7266, f(x) = 0.0000
          12'hA24: exp_out = 32'h00004448; // x = -11.7188, f(x) = 0.0000
          12'hA25: exp_out = 32'h000044D1; // x = -11.7109, f(x) = 0.0000
          12'hA26: exp_out = 32'h0000455B; // x = -11.7031, f(x) = 0.0000
          12'hA27: exp_out = 32'h000045E7; // x = -11.6953, f(x) = 0.0000
          12'hA28: exp_out = 32'h00004673; // x = -11.6875, f(x) = 0.0000
          12'hA29: exp_out = 32'h00004700; // x = -11.6797, f(x) = 0.0000
          12'hA2A: exp_out = 32'h0000478F; // x = -11.6719, f(x) = 0.0000
          12'hA2B: exp_out = 32'h0000481F; // x = -11.6641, f(x) = 0.0000
          12'hA2C: exp_out = 32'h000048AF; // x = -11.6562, f(x) = 0.0000
          12'hA2D: exp_out = 32'h00004941; // x = -11.6484, f(x) = 0.0000
          12'hA2E: exp_out = 32'h000049D4; // x = -11.6406, f(x) = 0.0000
          12'hA2F: exp_out = 32'h00004A69; // x = -11.6328, f(x) = 0.0000
          12'hA30: exp_out = 32'h00004AFE; // x = -11.6250, f(x) = 0.0000
          12'hA31: exp_out = 32'h00004B95; // x = -11.6172, f(x) = 0.0000
          12'hA32: exp_out = 32'h00004C2C; // x = -11.6094, f(x) = 0.0000
          12'hA33: exp_out = 32'h00004CC5; // x = -11.6016, f(x) = 0.0000
          12'hA34: exp_out = 32'h00004D5F; // x = -11.5938, f(x) = 0.0000
          12'hA35: exp_out = 32'h00004DFB; // x = -11.5859, f(x) = 0.0000
          12'hA36: exp_out = 32'h00004E97; // x = -11.5781, f(x) = 0.0000
          12'hA37: exp_out = 32'h00004F35; // x = -11.5703, f(x) = 0.0000
          12'hA38: exp_out = 32'h00004FD4; // x = -11.5625, f(x) = 0.0000
          12'hA39: exp_out = 32'h00005074; // x = -11.5547, f(x) = 0.0000
          12'hA3A: exp_out = 32'h00005116; // x = -11.5469, f(x) = 0.0000
          12'hA3B: exp_out = 32'h000051B9; // x = -11.5391, f(x) = 0.0000
          12'hA3C: exp_out = 32'h0000525D; // x = -11.5312, f(x) = 0.0000
          12'hA3D: exp_out = 32'h00005302; // x = -11.5234, f(x) = 0.0000
          12'hA3E: exp_out = 32'h000053A9; // x = -11.5156, f(x) = 0.0000
          12'hA3F: exp_out = 32'h00005451; // x = -11.5078, f(x) = 0.0000
          12'hA40: exp_out = 32'h000054FA; // x = -11.5000, f(x) = 0.0000
          12'hA41: exp_out = 32'h000055A5; // x = -11.4922, f(x) = 0.0000
          12'hA42: exp_out = 32'h00005651; // x = -11.4844, f(x) = 0.0000
          12'hA43: exp_out = 32'h000056FE; // x = -11.4766, f(x) = 0.0000
          12'hA44: exp_out = 32'h000057AD; // x = -11.4688, f(x) = 0.0000
          12'hA45: exp_out = 32'h0000585D; // x = -11.4609, f(x) = 0.0000
          12'hA46: exp_out = 32'h0000590E; // x = -11.4531, f(x) = 0.0000
          12'hA47: exp_out = 32'h000059C1; // x = -11.4453, f(x) = 0.0000
          12'hA48: exp_out = 32'h00005A75; // x = -11.4375, f(x) = 0.0000
          12'hA49: exp_out = 32'h00005B2B; // x = -11.4297, f(x) = 0.0000
          12'hA4A: exp_out = 32'h00005BE2; // x = -11.4219, f(x) = 0.0000
          12'hA4B: exp_out = 32'h00005C9A; // x = -11.4141, f(x) = 0.0000
          12'hA4C: exp_out = 32'h00005D54; // x = -11.4062, f(x) = 0.0000
          12'hA4D: exp_out = 32'h00005E10; // x = -11.3984, f(x) = 0.0000
          12'hA4E: exp_out = 32'h00005ECD; // x = -11.3906, f(x) = 0.0000
          12'hA4F: exp_out = 32'h00005F8B; // x = -11.3828, f(x) = 0.0000
          12'hA50: exp_out = 32'h0000604B; // x = -11.3750, f(x) = 0.0000
          12'hA51: exp_out = 32'h0000610C; // x = -11.3672, f(x) = 0.0000
          12'hA52: exp_out = 32'h000061CF; // x = -11.3594, f(x) = 0.0000
          12'hA53: exp_out = 32'h00006293; // x = -11.3516, f(x) = 0.0000
          12'hA54: exp_out = 32'h00006359; // x = -11.3438, f(x) = 0.0000
          12'hA55: exp_out = 32'h00006421; // x = -11.3359, f(x) = 0.0000
          12'hA56: exp_out = 32'h000064EA; // x = -11.3281, f(x) = 0.0000
          12'hA57: exp_out = 32'h000065B4; // x = -11.3203, f(x) = 0.0000
          12'hA58: exp_out = 32'h00006681; // x = -11.3125, f(x) = 0.0000
          12'hA59: exp_out = 32'h0000674E; // x = -11.3047, f(x) = 0.0000
          12'hA5A: exp_out = 32'h0000681E; // x = -11.2969, f(x) = 0.0000
          12'hA5B: exp_out = 32'h000068EF; // x = -11.2891, f(x) = 0.0000
          12'hA5C: exp_out = 32'h000069C2; // x = -11.2812, f(x) = 0.0000
          12'hA5D: exp_out = 32'h00006A96; // x = -11.2734, f(x) = 0.0000
          12'hA5E: exp_out = 32'h00006B6C; // x = -11.2656, f(x) = 0.0000
          12'hA5F: exp_out = 32'h00006C44; // x = -11.2578, f(x) = 0.0000
          12'hA60: exp_out = 32'h00006D1D; // x = -11.2500, f(x) = 0.0000
          12'hA61: exp_out = 32'h00006DF8; // x = -11.2422, f(x) = 0.0000
          12'hA62: exp_out = 32'h00006ED5; // x = -11.2344, f(x) = 0.0000
          12'hA63: exp_out = 32'h00006FB3; // x = -11.2266, f(x) = 0.0000
          12'hA64: exp_out = 32'h00007094; // x = -11.2188, f(x) = 0.0000
          12'hA65: exp_out = 32'h00007176; // x = -11.2109, f(x) = 0.0000
          12'hA66: exp_out = 32'h00007259; // x = -11.2031, f(x) = 0.0000
          12'hA67: exp_out = 32'h0000733F; // x = -11.1953, f(x) = 0.0000
          12'hA68: exp_out = 32'h00007426; // x = -11.1875, f(x) = 0.0000
          12'hA69: exp_out = 32'h00007510; // x = -11.1797, f(x) = 0.0000
          12'hA6A: exp_out = 32'h000075FB; // x = -11.1719, f(x) = 0.0000
          12'hA6B: exp_out = 32'h000076E8; // x = -11.1641, f(x) = 0.0000
          12'hA6C: exp_out = 32'h000077D6; // x = -11.1562, f(x) = 0.0000
          12'hA6D: exp_out = 32'h000078C7; // x = -11.1484, f(x) = 0.0000
          12'hA6E: exp_out = 32'h000079B9; // x = -11.1406, f(x) = 0.0000
          12'hA6F: exp_out = 32'h00007AAE; // x = -11.1328, f(x) = 0.0000
          12'hA70: exp_out = 32'h00007BA4; // x = -11.1250, f(x) = 0.0000
          12'hA71: exp_out = 32'h00007C9C; // x = -11.1172, f(x) = 0.0000
          12'hA72: exp_out = 32'h00007D97; // x = -11.1094, f(x) = 0.0000
          12'hA73: exp_out = 32'h00007E93; // x = -11.1016, f(x) = 0.0000
          12'hA74: exp_out = 32'h00007F91; // x = -11.0938, f(x) = 0.0000
          12'hA75: exp_out = 32'h00008091; // x = -11.0859, f(x) = 0.0000
          12'hA76: exp_out = 32'h00008193; // x = -11.0781, f(x) = 0.0000
          12'hA77: exp_out = 32'h00008297; // x = -11.0703, f(x) = 0.0000
          12'hA78: exp_out = 32'h0000839E; // x = -11.0625, f(x) = 0.0000
          12'hA79: exp_out = 32'h000084A6; // x = -11.0547, f(x) = 0.0000
          12'hA7A: exp_out = 32'h000085B0; // x = -11.0469, f(x) = 0.0000
          12'hA7B: exp_out = 32'h000086BD; // x = -11.0391, f(x) = 0.0000
          12'hA7C: exp_out = 32'h000087CB; // x = -11.0312, f(x) = 0.0000
          12'hA7D: exp_out = 32'h000088DC; // x = -11.0234, f(x) = 0.0000
          12'hA7E: exp_out = 32'h000089EF; // x = -11.0156, f(x) = 0.0000
          12'hA7F: exp_out = 32'h00008B04; // x = -11.0078, f(x) = 0.0000
          12'hA80: exp_out = 32'h00008C1B; // x = -11.0000, f(x) = 0.0000
          12'hA81: exp_out = 32'h00008D34; // x = -10.9922, f(x) = 0.0000
          12'hA82: exp_out = 32'h00008E4F; // x = -10.9844, f(x) = 0.0000
          12'hA83: exp_out = 32'h00008F6D; // x = -10.9766, f(x) = 0.0000
          12'hA84: exp_out = 32'h0000908D; // x = -10.9688, f(x) = 0.0000
          12'hA85: exp_out = 32'h000091AF; // x = -10.9609, f(x) = 0.0000
          12'hA86: exp_out = 32'h000092D4; // x = -10.9531, f(x) = 0.0000
          12'hA87: exp_out = 32'h000093FB; // x = -10.9453, f(x) = 0.0000
          12'hA88: exp_out = 32'h00009524; // x = -10.9375, f(x) = 0.0000
          12'hA89: exp_out = 32'h0000964F; // x = -10.9297, f(x) = 0.0000
          12'hA8A: exp_out = 32'h0000977D; // x = -10.9219, f(x) = 0.0000
          12'hA8B: exp_out = 32'h000098AD; // x = -10.9141, f(x) = 0.0000
          12'hA8C: exp_out = 32'h000099E0; // x = -10.9062, f(x) = 0.0000
          12'hA8D: exp_out = 32'h00009B15; // x = -10.8984, f(x) = 0.0000
          12'hA8E: exp_out = 32'h00009C4C; // x = -10.8906, f(x) = 0.0000
          12'hA8F: exp_out = 32'h00009D86; // x = -10.8828, f(x) = 0.0000
          12'hA90: exp_out = 32'h00009EC2; // x = -10.8750, f(x) = 0.0000
          12'hA91: exp_out = 32'h0000A001; // x = -10.8672, f(x) = 0.0000
          12'hA92: exp_out = 32'h0000A142; // x = -10.8594, f(x) = 0.0000
          12'hA93: exp_out = 32'h0000A286; // x = -10.8516, f(x) = 0.0000
          12'hA94: exp_out = 32'h0000A3CC; // x = -10.8438, f(x) = 0.0000
          12'hA95: exp_out = 32'h0000A515; // x = -10.8359, f(x) = 0.0000
          12'hA96: exp_out = 32'h0000A661; // x = -10.8281, f(x) = 0.0000
          12'hA97: exp_out = 32'h0000A7AF; // x = -10.8203, f(x) = 0.0000
          12'hA98: exp_out = 32'h0000A8FF; // x = -10.8125, f(x) = 0.0000
          12'hA99: exp_out = 32'h0000AA53; // x = -10.8047, f(x) = 0.0000
          12'hA9A: exp_out = 32'h0000ABA9; // x = -10.7969, f(x) = 0.0000
          12'hA9B: exp_out = 32'h0000AD01; // x = -10.7891, f(x) = 0.0000
          12'hA9C: exp_out = 32'h0000AE5D; // x = -10.7812, f(x) = 0.0000
          12'hA9D: exp_out = 32'h0000AFBB; // x = -10.7734, f(x) = 0.0000
          12'hA9E: exp_out = 32'h0000B11C; // x = -10.7656, f(x) = 0.0000
          12'hA9F: exp_out = 32'h0000B27F; // x = -10.7578, f(x) = 0.0000
          12'hAA0: exp_out = 32'h0000B3E6; // x = -10.7500, f(x) = 0.0000
          12'hAA1: exp_out = 32'h0000B54F; // x = -10.7422, f(x) = 0.0000
          12'hAA2: exp_out = 32'h0000B6BB; // x = -10.7344, f(x) = 0.0000
          12'hAA3: exp_out = 32'h0000B82A; // x = -10.7266, f(x) = 0.0000
          12'hAA4: exp_out = 32'h0000B99C; // x = -10.7188, f(x) = 0.0000
          12'hAA5: exp_out = 32'h0000BB10; // x = -10.7109, f(x) = 0.0000
          12'hAA6: exp_out = 32'h0000BC88; // x = -10.7031, f(x) = 0.0000
          12'hAA7: exp_out = 32'h0000BE02; // x = -10.6953, f(x) = 0.0000
          12'hAA8: exp_out = 32'h0000BF80; // x = -10.6875, f(x) = 0.0000
          12'hAA9: exp_out = 32'h0000C100; // x = -10.6797, f(x) = 0.0000
          12'hAAA: exp_out = 32'h0000C284; // x = -10.6719, f(x) = 0.0000
          12'hAAB: exp_out = 32'h0000C40A; // x = -10.6641, f(x) = 0.0000
          12'hAAC: exp_out = 32'h0000C594; // x = -10.6562, f(x) = 0.0000
          12'hAAD: exp_out = 32'h0000C721; // x = -10.6484, f(x) = 0.0000
          12'hAAE: exp_out = 32'h0000C8B1; // x = -10.6406, f(x) = 0.0000
          12'hAAF: exp_out = 32'h0000CA44; // x = -10.6328, f(x) = 0.0000
          12'hAB0: exp_out = 32'h0000CBDA; // x = -10.6250, f(x) = 0.0000
          12'hAB1: exp_out = 32'h0000CD73; // x = -10.6172, f(x) = 0.0000
          12'hAB2: exp_out = 32'h0000CF0F; // x = -10.6094, f(x) = 0.0000
          12'hAB3: exp_out = 32'h0000D0AF; // x = -10.6016, f(x) = 0.0000
          12'hAB4: exp_out = 32'h0000D252; // x = -10.5938, f(x) = 0.0000
          12'hAB5: exp_out = 32'h0000D3F8; // x = -10.5859, f(x) = 0.0000
          12'hAB6: exp_out = 32'h0000D5A2; // x = -10.5781, f(x) = 0.0000
          12'hAB7: exp_out = 32'h0000D74F; // x = -10.5703, f(x) = 0.0000
          12'hAB8: exp_out = 32'h0000D8FF; // x = -10.5625, f(x) = 0.0000
          12'hAB9: exp_out = 32'h0000DAB3; // x = -10.5547, f(x) = 0.0000
          12'hABA: exp_out = 32'h0000DC6A; // x = -10.5469, f(x) = 0.0000
          12'hABB: exp_out = 32'h0000DE25; // x = -10.5391, f(x) = 0.0000
          12'hABC: exp_out = 32'h0000DFE3; // x = -10.5312, f(x) = 0.0000
          12'hABD: exp_out = 32'h0000E1A4; // x = -10.5234, f(x) = 0.0000
          12'hABE: exp_out = 32'h0000E369; // x = -10.5156, f(x) = 0.0000
          12'hABF: exp_out = 32'h0000E532; // x = -10.5078, f(x) = 0.0000
          12'hAC0: exp_out = 32'h0000E6FE; // x = -10.5000, f(x) = 0.0000
          12'hAC1: exp_out = 32'h0000E8CE; // x = -10.4922, f(x) = 0.0000
          12'hAC2: exp_out = 32'h0000EAA1; // x = -10.4844, f(x) = 0.0000
          12'hAC3: exp_out = 32'h0000EC78; // x = -10.4766, f(x) = 0.0000
          12'hAC4: exp_out = 32'h0000EE53; // x = -10.4688, f(x) = 0.0000
          12'hAC5: exp_out = 32'h0000F032; // x = -10.4609, f(x) = 0.0000
          12'hAC6: exp_out = 32'h0000F214; // x = -10.4531, f(x) = 0.0000
          12'hAC7: exp_out = 32'h0000F3FA; // x = -10.4453, f(x) = 0.0000
          12'hAC8: exp_out = 32'h0000F5E4; // x = -10.4375, f(x) = 0.0000
          12'hAC9: exp_out = 32'h0000F7D2; // x = -10.4297, f(x) = 0.0000
          12'hACA: exp_out = 32'h0000F9C3; // x = -10.4219, f(x) = 0.0000
          12'hACB: exp_out = 32'h0000FBB9; // x = -10.4141, f(x) = 0.0000
          12'hACC: exp_out = 32'h0000FDB2; // x = -10.4062, f(x) = 0.0000
          12'hACD: exp_out = 32'h0000FFAF; // x = -10.3984, f(x) = 0.0000
          12'hACE: exp_out = 32'h000101B1; // x = -10.3906, f(x) = 0.0000
          12'hACF: exp_out = 32'h000103B6; // x = -10.3828, f(x) = 0.0000
          12'hAD0: exp_out = 32'h000105C0; // x = -10.3750, f(x) = 0.0000
          12'hAD1: exp_out = 32'h000107CD; // x = -10.3672, f(x) = 0.0000
          12'hAD2: exp_out = 32'h000109DF; // x = -10.3594, f(x) = 0.0000
          12'hAD3: exp_out = 32'h00010BF5; // x = -10.3516, f(x) = 0.0000
          12'hAD4: exp_out = 32'h00010E0F; // x = -10.3438, f(x) = 0.0000
          12'hAD5: exp_out = 32'h0001102D; // x = -10.3359, f(x) = 0.0000
          12'hAD6: exp_out = 32'h0001124F; // x = -10.3281, f(x) = 0.0000
          12'hAD7: exp_out = 32'h00011476; // x = -10.3203, f(x) = 0.0000
          12'hAD8: exp_out = 32'h000116A1; // x = -10.3125, f(x) = 0.0000
          12'hAD9: exp_out = 32'h000118D1; // x = -10.3047, f(x) = 0.0000
          12'hADA: exp_out = 32'h00011B05; // x = -10.2969, f(x) = 0.0000
          12'hADB: exp_out = 32'h00011D3D; // x = -10.2891, f(x) = 0.0000
          12'hADC: exp_out = 32'h00011F7A; // x = -10.2812, f(x) = 0.0000
          12'hADD: exp_out = 32'h000121BB; // x = -10.2734, f(x) = 0.0000
          12'hADE: exp_out = 32'h00012400; // x = -10.2656, f(x) = 0.0000
          12'hADF: exp_out = 32'h0001264B; // x = -10.2578, f(x) = 0.0000
          12'hAE0: exp_out = 32'h0001289A; // x = -10.2500, f(x) = 0.0000
          12'hAE1: exp_out = 32'h00012AED; // x = -10.2422, f(x) = 0.0000
          12'hAE2: exp_out = 32'h00012D45; // x = -10.2344, f(x) = 0.0000
          12'hAE3: exp_out = 32'h00012FA2; // x = -10.2266, f(x) = 0.0000
          12'hAE4: exp_out = 32'h00013204; // x = -10.2188, f(x) = 0.0000
          12'hAE5: exp_out = 32'h0001346A; // x = -10.2109, f(x) = 0.0000
          12'hAE6: exp_out = 32'h000136D6; // x = -10.2031, f(x) = 0.0000
          12'hAE7: exp_out = 32'h00013946; // x = -10.1953, f(x) = 0.0000
          12'hAE8: exp_out = 32'h00013BBB; // x = -10.1875, f(x) = 0.0000
          12'hAE9: exp_out = 32'h00013E35; // x = -10.1797, f(x) = 0.0000
          12'hAEA: exp_out = 32'h000140B4; // x = -10.1719, f(x) = 0.0000
          12'hAEB: exp_out = 32'h00014337; // x = -10.1641, f(x) = 0.0000
          12'hAEC: exp_out = 32'h000145C0; // x = -10.1562, f(x) = 0.0000
          12'hAED: exp_out = 32'h0001484E; // x = -10.1484, f(x) = 0.0000
          12'hAEE: exp_out = 32'h00014AE2; // x = -10.1406, f(x) = 0.0000
          12'hAEF: exp_out = 32'h00014D7A; // x = -10.1328, f(x) = 0.0000
          12'hAF0: exp_out = 32'h00015018; // x = -10.1250, f(x) = 0.0000
          12'hAF1: exp_out = 32'h000152BA; // x = -10.1172, f(x) = 0.0000
          12'hAF2: exp_out = 32'h00015562; // x = -10.1094, f(x) = 0.0000
          12'hAF3: exp_out = 32'h00015810; // x = -10.1016, f(x) = 0.0000
          12'hAF4: exp_out = 32'h00015AC3; // x = -10.0938, f(x) = 0.0000
          12'hAF5: exp_out = 32'h00015D7B; // x = -10.0859, f(x) = 0.0000
          12'hAF6: exp_out = 32'h00016039; // x = -10.0781, f(x) = 0.0000
          12'hAF7: exp_out = 32'h000162FC; // x = -10.0703, f(x) = 0.0000
          12'hAF8: exp_out = 32'h000165C5; // x = -10.0625, f(x) = 0.0000
          12'hAF9: exp_out = 32'h00016893; // x = -10.0547, f(x) = 0.0000
          12'hAFA: exp_out = 32'h00016B67; // x = -10.0469, f(x) = 0.0000
          12'hAFB: exp_out = 32'h00016E41; // x = -10.0391, f(x) = 0.0000
          12'hAFC: exp_out = 32'h00017120; // x = -10.0312, f(x) = 0.0000
          12'hAFD: exp_out = 32'h00017405; // x = -10.0234, f(x) = 0.0000
          12'hAFE: exp_out = 32'h000176F0; // x = -10.0156, f(x) = 0.0000
          12'hAFF: exp_out = 32'h000179E1; // x = -10.0078, f(x) = 0.0000
          12'hB00: exp_out = 32'h00017CD8; // x = -10.0000, f(x) = 0.0000
          12'hB01: exp_out = 32'h00017FD4; // x = -9.9922, f(x) = 0.0000
          12'hB02: exp_out = 32'h000182D7; // x = -9.9844, f(x) = 0.0000
          12'hB03: exp_out = 32'h000185E0; // x = -9.9766, f(x) = 0.0000
          12'hB04: exp_out = 32'h000188EE; // x = -9.9688, f(x) = 0.0000
          12'hB05: exp_out = 32'h00018C03; // x = -9.9609, f(x) = 0.0000
          12'hB06: exp_out = 32'h00018F1F; // x = -9.9531, f(x) = 0.0000
          12'hB07: exp_out = 32'h00019240; // x = -9.9453, f(x) = 0.0000
          12'hB08: exp_out = 32'h00019568; // x = -9.9375, f(x) = 0.0000
          12'hB09: exp_out = 32'h00019896; // x = -9.9297, f(x) = 0.0000
          12'hB0A: exp_out = 32'h00019BCA; // x = -9.9219, f(x) = 0.0000
          12'hB0B: exp_out = 32'h00019F05; // x = -9.9141, f(x) = 0.0000
          12'hB0C: exp_out = 32'h0001A246; // x = -9.9062, f(x) = 0.0000
          12'hB0D: exp_out = 32'h0001A58E; // x = -9.8984, f(x) = 0.0001
          12'hB0E: exp_out = 32'h0001A8DC; // x = -9.8906, f(x) = 0.0001
          12'hB0F: exp_out = 32'h0001AC31; // x = -9.8828, f(x) = 0.0001
          12'hB10: exp_out = 32'h0001AF8D; // x = -9.8750, f(x) = 0.0001
          12'hB11: exp_out = 32'h0001B2EF; // x = -9.8672, f(x) = 0.0001
          12'hB12: exp_out = 32'h0001B659; // x = -9.8594, f(x) = 0.0001
          12'hB13: exp_out = 32'h0001B9C9; // x = -9.8516, f(x) = 0.0001
          12'hB14: exp_out = 32'h0001BD40; // x = -9.8438, f(x) = 0.0001
          12'hB15: exp_out = 32'h0001C0BE; // x = -9.8359, f(x) = 0.0001
          12'hB16: exp_out = 32'h0001C443; // x = -9.8281, f(x) = 0.0001
          12'hB17: exp_out = 32'h0001C7CF; // x = -9.8203, f(x) = 0.0001
          12'hB18: exp_out = 32'h0001CB62; // x = -9.8125, f(x) = 0.0001
          12'hB19: exp_out = 32'h0001CEFD; // x = -9.8047, f(x) = 0.0001
          12'hB1A: exp_out = 32'h0001D29E; // x = -9.7969, f(x) = 0.0001
          12'hB1B: exp_out = 32'h0001D647; // x = -9.7891, f(x) = 0.0001
          12'hB1C: exp_out = 32'h0001D9F7; // x = -9.7812, f(x) = 0.0001
          12'hB1D: exp_out = 32'h0001DDAF; // x = -9.7734, f(x) = 0.0001
          12'hB1E: exp_out = 32'h0001E16E; // x = -9.7656, f(x) = 0.0001
          12'hB1F: exp_out = 32'h0001E535; // x = -9.7578, f(x) = 0.0001
          12'hB20: exp_out = 32'h0001E903; // x = -9.7500, f(x) = 0.0001
          12'hB21: exp_out = 32'h0001ECD9; // x = -9.7422, f(x) = 0.0001
          12'hB22: exp_out = 32'h0001F0B6; // x = -9.7344, f(x) = 0.0001
          12'hB23: exp_out = 32'h0001F49C; // x = -9.7266, f(x) = 0.0001
          12'hB24: exp_out = 32'h0001F889; // x = -9.7188, f(x) = 0.0001
          12'hB25: exp_out = 32'h0001FC7E; // x = -9.7109, f(x) = 0.0001
          12'hB26: exp_out = 32'h0002007B; // x = -9.7031, f(x) = 0.0001
          12'hB27: exp_out = 32'h00020480; // x = -9.6953, f(x) = 0.0001
          12'hB28: exp_out = 32'h0002088D; // x = -9.6875, f(x) = 0.0001
          12'hB29: exp_out = 32'h00020CA2; // x = -9.6797, f(x) = 0.0001
          12'hB2A: exp_out = 32'h000210BF; // x = -9.6719, f(x) = 0.0001
          12'hB2B: exp_out = 32'h000214E5; // x = -9.6641, f(x) = 0.0001
          12'hB2C: exp_out = 32'h00021913; // x = -9.6562, f(x) = 0.0001
          12'hB2D: exp_out = 32'h00021D49; // x = -9.6484, f(x) = 0.0001
          12'hB2E: exp_out = 32'h00022188; // x = -9.6406, f(x) = 0.0001
          12'hB2F: exp_out = 32'h000225CF; // x = -9.6328, f(x) = 0.0001
          12'hB30: exp_out = 32'h00022A1F; // x = -9.6250, f(x) = 0.0001
          12'hB31: exp_out = 32'h00022E78; // x = -9.6172, f(x) = 0.0001
          12'hB32: exp_out = 32'h000232D9; // x = -9.6094, f(x) = 0.0001
          12'hB33: exp_out = 32'h00023743; // x = -9.6016, f(x) = 0.0001
          12'hB34: exp_out = 32'h00023BB6; // x = -9.5938, f(x) = 0.0001
          12'hB35: exp_out = 32'h00024032; // x = -9.5859, f(x) = 0.0001
          12'hB36: exp_out = 32'h000244B7; // x = -9.5781, f(x) = 0.0001
          12'hB37: exp_out = 32'h00024945; // x = -9.5703, f(x) = 0.0001
          12'hB38: exp_out = 32'h00024DDC; // x = -9.5625, f(x) = 0.0001
          12'hB39: exp_out = 32'h0002527C; // x = -9.5547, f(x) = 0.0001
          12'hB3A: exp_out = 32'h00025726; // x = -9.5469, f(x) = 0.0001
          12'hB3B: exp_out = 32'h00025BD9; // x = -9.5391, f(x) = 0.0001
          12'hB3C: exp_out = 32'h00026096; // x = -9.5312, f(x) = 0.0001
          12'hB3D: exp_out = 32'h0002655B; // x = -9.5234, f(x) = 0.0001
          12'hB3E: exp_out = 32'h00026A2B; // x = -9.5156, f(x) = 0.0001
          12'hB3F: exp_out = 32'h00026F04; // x = -9.5078, f(x) = 0.0001
          12'hB40: exp_out = 32'h000273E7; // x = -9.5000, f(x) = 0.0001
          12'hB41: exp_out = 32'h000278D4; // x = -9.4922, f(x) = 0.0001
          12'hB42: exp_out = 32'h00027DCA; // x = -9.4844, f(x) = 0.0001
          12'hB43: exp_out = 32'h000282CB; // x = -9.4766, f(x) = 0.0001
          12'hB44: exp_out = 32'h000287D6; // x = -9.4688, f(x) = 0.0001
          12'hB45: exp_out = 32'h00028CEA; // x = -9.4609, f(x) = 0.0001
          12'hB46: exp_out = 32'h00029209; // x = -9.4531, f(x) = 0.0001
          12'hB47: exp_out = 32'h00029733; // x = -9.4453, f(x) = 0.0001
          12'hB48: exp_out = 32'h00029C66; // x = -9.4375, f(x) = 0.0001
          12'hB49: exp_out = 32'h0002A1A4; // x = -9.4297, f(x) = 0.0001
          12'hB4A: exp_out = 32'h0002A6ED; // x = -9.4219, f(x) = 0.0001
          12'hB4B: exp_out = 32'h0002AC40; // x = -9.4141, f(x) = 0.0001
          12'hB4C: exp_out = 32'h0002B19E; // x = -9.4062, f(x) = 0.0001
          12'hB4D: exp_out = 32'h0002B706; // x = -9.3984, f(x) = 0.0001
          12'hB4E: exp_out = 32'h0002BC7A; // x = -9.3906, f(x) = 0.0001
          12'hB4F: exp_out = 32'h0002C1F8; // x = -9.3828, f(x) = 0.0001
          12'hB50: exp_out = 32'h0002C782; // x = -9.3750, f(x) = 0.0001
          12'hB51: exp_out = 32'h0002CD16; // x = -9.3672, f(x) = 0.0001
          12'hB52: exp_out = 32'h0002D2B6; // x = -9.3594, f(x) = 0.0001
          12'hB53: exp_out = 32'h0002D861; // x = -9.3516, f(x) = 0.0001
          12'hB54: exp_out = 32'h0002DE18; // x = -9.3438, f(x) = 0.0001
          12'hB55: exp_out = 32'h0002E3DA; // x = -9.3359, f(x) = 0.0001
          12'hB56: exp_out = 32'h0002E9A7; // x = -9.3281, f(x) = 0.0001
          12'hB57: exp_out = 32'h0002EF80; // x = -9.3203, f(x) = 0.0001
          12'hB58: exp_out = 32'h0002F565; // x = -9.3125, f(x) = 0.0001
          12'hB59: exp_out = 32'h0002FB56; // x = -9.3047, f(x) = 0.0001
          12'hB5A: exp_out = 32'h00030153; // x = -9.2969, f(x) = 0.0001
          12'hB5B: exp_out = 32'h0003075B; // x = -9.2891, f(x) = 0.0001
          12'hB5C: exp_out = 32'h00030D70; // x = -9.2812, f(x) = 0.0001
          12'hB5D: exp_out = 32'h00031391; // x = -9.2734, f(x) = 0.0001
          12'hB5E: exp_out = 32'h000319BE; // x = -9.2656, f(x) = 0.0001
          12'hB5F: exp_out = 32'h00031FF8; // x = -9.2578, f(x) = 0.0001
          12'hB60: exp_out = 32'h0003263E; // x = -9.2500, f(x) = 0.0001
          12'hB61: exp_out = 32'h00032C91; // x = -9.2422, f(x) = 0.0001
          12'hB62: exp_out = 32'h000332F0; // x = -9.2344, f(x) = 0.0001
          12'hB63: exp_out = 32'h0003395D; // x = -9.2266, f(x) = 0.0001
          12'hB64: exp_out = 32'h00033FD6; // x = -9.2188, f(x) = 0.0001
          12'hB65: exp_out = 32'h0003465C; // x = -9.2109, f(x) = 0.0001
          12'hB66: exp_out = 32'h00034CEF; // x = -9.2031, f(x) = 0.0001
          12'hB67: exp_out = 32'h00035390; // x = -9.1953, f(x) = 0.0001
          12'hB68: exp_out = 32'h00035A3E; // x = -9.1875, f(x) = 0.0001
          12'hB69: exp_out = 32'h000360F9; // x = -9.1797, f(x) = 0.0001
          12'hB6A: exp_out = 32'h000367C2; // x = -9.1719, f(x) = 0.0001
          12'hB6B: exp_out = 32'h00036E98; // x = -9.1641, f(x) = 0.0001
          12'hB6C: exp_out = 32'h0003757C; // x = -9.1562, f(x) = 0.0001
          12'hB6D: exp_out = 32'h00037C6E; // x = -9.1484, f(x) = 0.0001
          12'hB6E: exp_out = 32'h0003836E; // x = -9.1406, f(x) = 0.0001
          12'hB6F: exp_out = 32'h00038A7C; // x = -9.1328, f(x) = 0.0001
          12'hB70: exp_out = 32'h00039198; // x = -9.1250, f(x) = 0.0001
          12'hB71: exp_out = 32'h000398C2; // x = -9.1172, f(x) = 0.0001
          12'hB72: exp_out = 32'h00039FFB; // x = -9.1094, f(x) = 0.0001
          12'hB73: exp_out = 32'h0003A742; // x = -9.1016, f(x) = 0.0001
          12'hB74: exp_out = 32'h0003AE98; // x = -9.0938, f(x) = 0.0001
          12'hB75: exp_out = 32'h0003B5FD; // x = -9.0859, f(x) = 0.0001
          12'hB76: exp_out = 32'h0003BD70; // x = -9.0781, f(x) = 0.0001
          12'hB77: exp_out = 32'h0003C4F2; // x = -9.0703, f(x) = 0.0001
          12'hB78: exp_out = 32'h0003CC84; // x = -9.0625, f(x) = 0.0001
          12'hB79: exp_out = 32'h0003D424; // x = -9.0547, f(x) = 0.0001
          12'hB7A: exp_out = 32'h0003DBD4; // x = -9.0469, f(x) = 0.0001
          12'hB7B: exp_out = 32'h0003E394; // x = -9.0391, f(x) = 0.0001
          12'hB7C: exp_out = 32'h0003EB63; // x = -9.0312, f(x) = 0.0001
          12'hB7D: exp_out = 32'h0003F341; // x = -9.0234, f(x) = 0.0001
          12'hB7E: exp_out = 32'h0003FB30; // x = -9.0156, f(x) = 0.0001
          12'hB7F: exp_out = 32'h0004032E; // x = -9.0078, f(x) = 0.0001
          12'hB80: exp_out = 32'h00040B3D; // x = -9.0000, f(x) = 0.0001
          12'hB81: exp_out = 32'h0004135B; // x = -8.9922, f(x) = 0.0001
          12'hB82: exp_out = 32'h00041B8A; // x = -8.9844, f(x) = 0.0001
          12'hB83: exp_out = 32'h000423C9; // x = -8.9766, f(x) = 0.0001
          12'hB84: exp_out = 32'h00042C19; // x = -8.9688, f(x) = 0.0001
          12'hB85: exp_out = 32'h0004347A; // x = -8.9609, f(x) = 0.0001
          12'hB86: exp_out = 32'h00043CEB; // x = -8.9531, f(x) = 0.0001
          12'hB87: exp_out = 32'h0004456D; // x = -8.9453, f(x) = 0.0001
          12'hB88: exp_out = 32'h00044E01; // x = -8.9375, f(x) = 0.0001
          12'hB89: exp_out = 32'h000456A6; // x = -8.9297, f(x) = 0.0001
          12'hB8A: exp_out = 32'h00045F5C; // x = -8.9219, f(x) = 0.0001
          12'hB8B: exp_out = 32'h00046823; // x = -8.9141, f(x) = 0.0001
          12'hB8C: exp_out = 32'h000470FC; // x = -8.9062, f(x) = 0.0001
          12'hB8D: exp_out = 32'h000479E7; // x = -8.8984, f(x) = 0.0001
          12'hB8E: exp_out = 32'h000482E4; // x = -8.8906, f(x) = 0.0001
          12'hB8F: exp_out = 32'h00048BF3; // x = -8.8828, f(x) = 0.0001
          12'hB90: exp_out = 32'h00049514; // x = -8.8750, f(x) = 0.0001
          12'hB91: exp_out = 32'h00049E47; // x = -8.8672, f(x) = 0.0001
          12'hB92: exp_out = 32'h0004A78D; // x = -8.8594, f(x) = 0.0001
          12'hB93: exp_out = 32'h0004B0E5; // x = -8.8516, f(x) = 0.0001
          12'hB94: exp_out = 32'h0004BA50; // x = -8.8438, f(x) = 0.0001
          12'hB95: exp_out = 32'h0004C3CF; // x = -8.8359, f(x) = 0.0001
          12'hB96: exp_out = 32'h0004CD60; // x = -8.8281, f(x) = 0.0001
          12'hB97: exp_out = 32'h0004D704; // x = -8.8203, f(x) = 0.0001
          12'hB98: exp_out = 32'h0004E0BC; // x = -8.8125, f(x) = 0.0001
          12'hB99: exp_out = 32'h0004EA87; // x = -8.8047, f(x) = 0.0002
          12'hB9A: exp_out = 32'h0004F466; // x = -8.7969, f(x) = 0.0002
          12'hB9B: exp_out = 32'h0004FE59; // x = -8.7891, f(x) = 0.0002
          12'hB9C: exp_out = 32'h0005085F; // x = -8.7812, f(x) = 0.0002
          12'hB9D: exp_out = 32'h0005127A; // x = -8.7734, f(x) = 0.0002
          12'hB9E: exp_out = 32'h00051CA9; // x = -8.7656, f(x) = 0.0002
          12'hB9F: exp_out = 32'h000526ED; // x = -8.7578, f(x) = 0.0002
          12'hBA0: exp_out = 32'h00053145; // x = -8.7500, f(x) = 0.0002
          12'hBA1: exp_out = 32'h00053BB2; // x = -8.7422, f(x) = 0.0002
          12'hBA2: exp_out = 32'h00054634; // x = -8.7344, f(x) = 0.0002
          12'hBA3: exp_out = 32'h000550CB; // x = -8.7266, f(x) = 0.0002
          12'hBA4: exp_out = 32'h00055B77; // x = -8.7188, f(x) = 0.0002
          12'hBA5: exp_out = 32'h00056639; // x = -8.7109, f(x) = 0.0002
          12'hBA6: exp_out = 32'h00057110; // x = -8.7031, f(x) = 0.0002
          12'hBA7: exp_out = 32'h00057BFD; // x = -8.6953, f(x) = 0.0002
          12'hBA8: exp_out = 32'h00058700; // x = -8.6875, f(x) = 0.0002
          12'hBA9: exp_out = 32'h00059219; // x = -8.6797, f(x) = 0.0002
          12'hBAA: exp_out = 32'h00059D49; // x = -8.6719, f(x) = 0.0002
          12'hBAB: exp_out = 32'h0005A88E; // x = -8.6641, f(x) = 0.0002
          12'hBAC: exp_out = 32'h0005B3EB; // x = -8.6562, f(x) = 0.0002
          12'hBAD: exp_out = 32'h0005BF5E; // x = -8.6484, f(x) = 0.0002
          12'hBAE: exp_out = 32'h0005CAE8; // x = -8.6406, f(x) = 0.0002
          12'hBAF: exp_out = 32'h0005D68A; // x = -8.6328, f(x) = 0.0002
          12'hBB0: exp_out = 32'h0005E243; // x = -8.6250, f(x) = 0.0002
          12'hBB1: exp_out = 32'h0005EE13; // x = -8.6172, f(x) = 0.0002
          12'hBB2: exp_out = 32'h0005F9FB; // x = -8.6094, f(x) = 0.0002
          12'hBB3: exp_out = 32'h000605FB; // x = -8.6016, f(x) = 0.0002
          12'hBB4: exp_out = 32'h00061213; // x = -8.5938, f(x) = 0.0002
          12'hBB5: exp_out = 32'h00061E43; // x = -8.5859, f(x) = 0.0002
          12'hBB6: exp_out = 32'h00062A8C; // x = -8.5781, f(x) = 0.0002
          12'hBB7: exp_out = 32'h000636EE; // x = -8.5703, f(x) = 0.0002
          12'hBB8: exp_out = 32'h00064368; // x = -8.5625, f(x) = 0.0002
          12'hBB9: exp_out = 32'h00064FFB; // x = -8.5547, f(x) = 0.0002
          12'hBBA: exp_out = 32'h00065CA8; // x = -8.5469, f(x) = 0.0002
          12'hBBB: exp_out = 32'h0006696E; // x = -8.5391, f(x) = 0.0002
          12'hBBC: exp_out = 32'h0006764E; // x = -8.5312, f(x) = 0.0002
          12'hBBD: exp_out = 32'h00068347; // x = -8.5234, f(x) = 0.0002
          12'hBBE: exp_out = 32'h0006905B; // x = -8.5156, f(x) = 0.0002
          12'hBBF: exp_out = 32'h00069D89; // x = -8.5078, f(x) = 0.0002
          12'hBC0: exp_out = 32'h0006AAD1; // x = -8.5000, f(x) = 0.0002
          12'hBC1: exp_out = 32'h0006B834; // x = -8.4922, f(x) = 0.0002
          12'hBC2: exp_out = 32'h0006C5B2; // x = -8.4844, f(x) = 0.0002
          12'hBC3: exp_out = 32'h0006D34B; // x = -8.4766, f(x) = 0.0002
          12'hBC4: exp_out = 32'h0006E0FF; // x = -8.4688, f(x) = 0.0002
          12'hBC5: exp_out = 32'h0006EECF; // x = -8.4609, f(x) = 0.0002
          12'hBC6: exp_out = 32'h0006FCBA; // x = -8.4531, f(x) = 0.0002
          12'hBC7: exp_out = 32'h00070AC2; // x = -8.4453, f(x) = 0.0002
          12'hBC8: exp_out = 32'h000718E6; // x = -8.4375, f(x) = 0.0002
          12'hBC9: exp_out = 32'h00072726; // x = -8.4297, f(x) = 0.0002
          12'hBCA: exp_out = 32'h00073582; // x = -8.4219, f(x) = 0.0002
          12'hBCB: exp_out = 32'h000743FC; // x = -8.4141, f(x) = 0.0002
          12'hBCC: exp_out = 32'h00075292; // x = -8.4062, f(x) = 0.0002
          12'hBCD: exp_out = 32'h00076146; // x = -8.3984, f(x) = 0.0002
          12'hBCE: exp_out = 32'h00077017; // x = -8.3906, f(x) = 0.0002
          12'hBCF: exp_out = 32'h00077F06; // x = -8.3828, f(x) = 0.0002
          12'hBD0: exp_out = 32'h00078E14; // x = -8.3750, f(x) = 0.0002
          12'hBD1: exp_out = 32'h00079D3F; // x = -8.3672, f(x) = 0.0002
          12'hBD2: exp_out = 32'h0007AC89; // x = -8.3594, f(x) = 0.0002
          12'hBD3: exp_out = 32'h0007BBF1; // x = -8.3516, f(x) = 0.0002
          12'hBD4: exp_out = 32'h0007CB78; // x = -8.3438, f(x) = 0.0002
          12'hBD5: exp_out = 32'h0007DB1F; // x = -8.3359, f(x) = 0.0002
          12'hBD6: exp_out = 32'h0007EAE5; // x = -8.3281, f(x) = 0.0002
          12'hBD7: exp_out = 32'h0007FACB; // x = -8.3203, f(x) = 0.0002
          12'hBD8: exp_out = 32'h00080AD0; // x = -8.3125, f(x) = 0.0002
          12'hBD9: exp_out = 32'h00081AF6; // x = -8.3047, f(x) = 0.0002
          12'hBDA: exp_out = 32'h00082B3C; // x = -8.2969, f(x) = 0.0002
          12'hBDB: exp_out = 32'h00083BA3; // x = -8.2891, f(x) = 0.0003
          12'hBDC: exp_out = 32'h00084C2B; // x = -8.2812, f(x) = 0.0003
          12'hBDD: exp_out = 32'h00085CD4; // x = -8.2734, f(x) = 0.0003
          12'hBDE: exp_out = 32'h00086D9E; // x = -8.2656, f(x) = 0.0003
          12'hBDF: exp_out = 32'h00087E8A; // x = -8.2578, f(x) = 0.0003
          12'hBE0: exp_out = 32'h00088F98; // x = -8.2500, f(x) = 0.0003
          12'hBE1: exp_out = 32'h0008A0C9; // x = -8.2422, f(x) = 0.0003
          12'hBE2: exp_out = 32'h0008B21C; // x = -8.2344, f(x) = 0.0003
          12'hBE3: exp_out = 32'h0008C391; // x = -8.2266, f(x) = 0.0003
          12'hBE4: exp_out = 32'h0008D52A; // x = -8.2188, f(x) = 0.0003
          12'hBE5: exp_out = 32'h0008E6E6; // x = -8.2109, f(x) = 0.0003
          12'hBE6: exp_out = 32'h0008F8C6; // x = -8.2031, f(x) = 0.0003
          12'hBE7: exp_out = 32'h00090AC9; // x = -8.1953, f(x) = 0.0003
          12'hBE8: exp_out = 32'h00091CF1; // x = -8.1875, f(x) = 0.0003
          12'hBE9: exp_out = 32'h00092F3D; // x = -8.1797, f(x) = 0.0003
          12'hBEA: exp_out = 32'h000941AE; // x = -8.1719, f(x) = 0.0003
          12'hBEB: exp_out = 32'h00095444; // x = -8.1641, f(x) = 0.0003
          12'hBEC: exp_out = 32'h000966FF; // x = -8.1562, f(x) = 0.0003
          12'hBED: exp_out = 32'h000979E0; // x = -8.1484, f(x) = 0.0003
          12'hBEE: exp_out = 32'h00098CE7; // x = -8.1406, f(x) = 0.0003
          12'hBEF: exp_out = 32'h0009A014; // x = -8.1328, f(x) = 0.0003
          12'hBF0: exp_out = 32'h0009B367; // x = -8.1250, f(x) = 0.0003
          12'hBF1: exp_out = 32'h0009C6E1; // x = -8.1172, f(x) = 0.0003
          12'hBF2: exp_out = 32'h0009DA83; // x = -8.1094, f(x) = 0.0003
          12'hBF3: exp_out = 32'h0009EE4C; // x = -8.1016, f(x) = 0.0003
          12'hBF4: exp_out = 32'h000A023C; // x = -8.0938, f(x) = 0.0003
          12'hBF5: exp_out = 32'h000A1655; // x = -8.0859, f(x) = 0.0003
          12'hBF6: exp_out = 32'h000A2A96; // x = -8.0781, f(x) = 0.0003
          12'hBF7: exp_out = 32'h000A3EFF; // x = -8.0703, f(x) = 0.0003
          12'hBF8: exp_out = 32'h000A5392; // x = -8.0625, f(x) = 0.0003
          12'hBF9: exp_out = 32'h000A684D; // x = -8.0547, f(x) = 0.0003
          12'hBFA: exp_out = 32'h000A7D33; // x = -8.0469, f(x) = 0.0003
          12'hBFB: exp_out = 32'h000A9242; // x = -8.0391, f(x) = 0.0003
          12'hBFC: exp_out = 32'h000AA77C; // x = -8.0312, f(x) = 0.0003
          12'hBFD: exp_out = 32'h000ABCE0; // x = -8.0234, f(x) = 0.0003
          12'hBFE: exp_out = 32'h000AD270; // x = -8.0156, f(x) = 0.0003
          12'hBFF: exp_out = 32'h000AE82A; // x = -8.0078, f(x) = 0.0003
          12'hC00: exp_out = 32'h000AFE11; // x = -8.0000, f(x) = 0.0003
          12'hC01: exp_out = 32'h000B1423; // x = -7.9922, f(x) = 0.0003
          12'hC02: exp_out = 32'h000B2A61; // x = -7.9844, f(x) = 0.0003
          12'hC03: exp_out = 32'h000B40CC; // x = -7.9766, f(x) = 0.0003
          12'hC04: exp_out = 32'h000B5764; // x = -7.9688, f(x) = 0.0003
          12'hC05: exp_out = 32'h000B6E2A; // x = -7.9609, f(x) = 0.0003
          12'hC06: exp_out = 32'h000B851D; // x = -7.9531, f(x) = 0.0004
          12'hC07: exp_out = 32'h000B9C3F; // x = -7.9453, f(x) = 0.0004
          12'hC08: exp_out = 32'h000BB38E; // x = -7.9375, f(x) = 0.0004
          12'hC09: exp_out = 32'h000BCB0D; // x = -7.9297, f(x) = 0.0004
          12'hC0A: exp_out = 32'h000BE2BB; // x = -7.9219, f(x) = 0.0004
          12'hC0B: exp_out = 32'h000BFA98; // x = -7.9141, f(x) = 0.0004
          12'hC0C: exp_out = 32'h000C12A5; // x = -7.9062, f(x) = 0.0004
          12'hC0D: exp_out = 32'h000C2AE3; // x = -7.8984, f(x) = 0.0004
          12'hC0E: exp_out = 32'h000C4351; // x = -7.8906, f(x) = 0.0004
          12'hC0F: exp_out = 32'h000C5BF0; // x = -7.8828, f(x) = 0.0004
          12'hC10: exp_out = 32'h000C74C1; // x = -7.8750, f(x) = 0.0004
          12'hC11: exp_out = 32'h000C8DC3; // x = -7.8672, f(x) = 0.0004
          12'hC12: exp_out = 32'h000CA6F8; // x = -7.8594, f(x) = 0.0004
          12'hC13: exp_out = 32'h000CC05F; // x = -7.8516, f(x) = 0.0004
          12'hC14: exp_out = 32'h000CD9FA; // x = -7.8438, f(x) = 0.0004
          12'hC15: exp_out = 32'h000CF3C7; // x = -7.8359, f(x) = 0.0004
          12'hC16: exp_out = 32'h000D0DC9; // x = -7.8281, f(x) = 0.0004
          12'hC17: exp_out = 32'h000D27FF; // x = -7.8203, f(x) = 0.0004
          12'hC18: exp_out = 32'h000D4269; // x = -7.8125, f(x) = 0.0004
          12'hC19: exp_out = 32'h000D5D08; // x = -7.8047, f(x) = 0.0004
          12'hC1A: exp_out = 32'h000D77DD; // x = -7.7969, f(x) = 0.0004
          12'hC1B: exp_out = 32'h000D92E8; // x = -7.7891, f(x) = 0.0004
          12'hC1C: exp_out = 32'h000DAE29; // x = -7.7812, f(x) = 0.0004
          12'hC1D: exp_out = 32'h000DC9A1; // x = -7.7734, f(x) = 0.0004
          12'hC1E: exp_out = 32'h000DE550; // x = -7.7656, f(x) = 0.0004
          12'hC1F: exp_out = 32'h000E0136; // x = -7.7578, f(x) = 0.0004
          12'hC20: exp_out = 32'h000E1D55; // x = -7.7500, f(x) = 0.0004
          12'hC21: exp_out = 32'h000E39AC; // x = -7.7422, f(x) = 0.0004
          12'hC22: exp_out = 32'h000E563B; // x = -7.7344, f(x) = 0.0004
          12'hC23: exp_out = 32'h000E7305; // x = -7.7266, f(x) = 0.0004
          12'hC24: exp_out = 32'h000E9008; // x = -7.7188, f(x) = 0.0004
          12'hC25: exp_out = 32'h000EAD45; // x = -7.7109, f(x) = 0.0004
          12'hC26: exp_out = 32'h000ECABD; // x = -7.7031, f(x) = 0.0005
          12'hC27: exp_out = 32'h000EE870; // x = -7.6953, f(x) = 0.0005
          12'hC28: exp_out = 32'h000F065F; // x = -7.6875, f(x) = 0.0005
          12'hC29: exp_out = 32'h000F248A; // x = -7.6797, f(x) = 0.0005
          12'hC2A: exp_out = 32'h000F42F1; // x = -7.6719, f(x) = 0.0005
          12'hC2B: exp_out = 32'h000F6196; // x = -7.6641, f(x) = 0.0005
          12'hC2C: exp_out = 32'h000F8078; // x = -7.6562, f(x) = 0.0005
          12'hC2D: exp_out = 32'h000F9F98; // x = -7.6484, f(x) = 0.0005
          12'hC2E: exp_out = 32'h000FBEF6; // x = -7.6406, f(x) = 0.0005
          12'hC2F: exp_out = 32'h000FDE94; // x = -7.6328, f(x) = 0.0005
          12'hC30: exp_out = 32'h000FFE71; // x = -7.6250, f(x) = 0.0005
          12'hC31: exp_out = 32'h00101E8E; // x = -7.6172, f(x) = 0.0005
          12'hC32: exp_out = 32'h00103EEB; // x = -7.6094, f(x) = 0.0005
          12'hC33: exp_out = 32'h00105F89; // x = -7.6016, f(x) = 0.0005
          12'hC34: exp_out = 32'h00108069; // x = -7.5938, f(x) = 0.0005
          12'hC35: exp_out = 32'h0010A18B; // x = -7.5859, f(x) = 0.0005
          12'hC36: exp_out = 32'h0010C2F0; // x = -7.5781, f(x) = 0.0005
          12'hC37: exp_out = 32'h0010E497; // x = -7.5703, f(x) = 0.0005
          12'hC38: exp_out = 32'h00110682; // x = -7.5625, f(x) = 0.0005
          12'hC39: exp_out = 32'h001128B1; // x = -7.5547, f(x) = 0.0005
          12'hC3A: exp_out = 32'h00114B25; // x = -7.5469, f(x) = 0.0005
          12'hC3B: exp_out = 32'h00116DDE; // x = -7.5391, f(x) = 0.0005
          12'hC3C: exp_out = 32'h001190DD; // x = -7.5312, f(x) = 0.0005
          12'hC3D: exp_out = 32'h0011B422; // x = -7.5234, f(x) = 0.0005
          12'hC3E: exp_out = 32'h0011D7AD; // x = -7.5156, f(x) = 0.0005
          12'hC3F: exp_out = 32'h0011FB81; // x = -7.5078, f(x) = 0.0005
          12'hC40: exp_out = 32'h00121F9C; // x = -7.5000, f(x) = 0.0006
          12'hC41: exp_out = 32'h001243FF; // x = -7.4922, f(x) = 0.0006
          12'hC42: exp_out = 32'h001268AC; // x = -7.4844, f(x) = 0.0006
          12'hC43: exp_out = 32'h00128DA2; // x = -7.4766, f(x) = 0.0006
          12'hC44: exp_out = 32'h0012B2E3; // x = -7.4688, f(x) = 0.0006
          12'hC45: exp_out = 32'h0012D86E; // x = -7.4609, f(x) = 0.0006
          12'hC46: exp_out = 32'h0012FE44; // x = -7.4531, f(x) = 0.0006
          12'hC47: exp_out = 32'h00132467; // x = -7.4453, f(x) = 0.0006
          12'hC48: exp_out = 32'h00134AD6; // x = -7.4375, f(x) = 0.0006
          12'hC49: exp_out = 32'h00137193; // x = -7.4297, f(x) = 0.0006
          12'hC4A: exp_out = 32'h0013989D; // x = -7.4219, f(x) = 0.0006
          12'hC4B: exp_out = 32'h0013BFF5; // x = -7.4141, f(x) = 0.0006
          12'hC4C: exp_out = 32'h0013E79D; // x = -7.4062, f(x) = 0.0006
          12'hC4D: exp_out = 32'h00140F94; // x = -7.3984, f(x) = 0.0006
          12'hC4E: exp_out = 32'h001437DB; // x = -7.3906, f(x) = 0.0006
          12'hC4F: exp_out = 32'h00146074; // x = -7.3828, f(x) = 0.0006
          12'hC50: exp_out = 32'h0014895D; // x = -7.3750, f(x) = 0.0006
          12'hC51: exp_out = 32'h0014B299; // x = -7.3672, f(x) = 0.0006
          12'hC52: exp_out = 32'h0014DC28; // x = -7.3594, f(x) = 0.0006
          12'hC53: exp_out = 32'h0015060A; // x = -7.3516, f(x) = 0.0006
          12'hC54: exp_out = 32'h00153040; // x = -7.3438, f(x) = 0.0006
          12'hC55: exp_out = 32'h00155ACB; // x = -7.3359, f(x) = 0.0007
          12'hC56: exp_out = 32'h001585AC; // x = -7.3281, f(x) = 0.0007
          12'hC57: exp_out = 32'h0015B0E2; // x = -7.3203, f(x) = 0.0007
          12'hC58: exp_out = 32'h0015DC6F; // x = -7.3125, f(x) = 0.0007
          12'hC59: exp_out = 32'h00160854; // x = -7.3047, f(x) = 0.0007
          12'hC5A: exp_out = 32'h00163491; // x = -7.2969, f(x) = 0.0007
          12'hC5B: exp_out = 32'h00166127; // x = -7.2891, f(x) = 0.0007
          12'hC5C: exp_out = 32'h00168E16; // x = -7.2812, f(x) = 0.0007
          12'hC5D: exp_out = 32'h0016BB5F; // x = -7.2734, f(x) = 0.0007
          12'hC5E: exp_out = 32'h0016E904; // x = -7.2656, f(x) = 0.0007
          12'hC5F: exp_out = 32'h00171704; // x = -7.2578, f(x) = 0.0007
          12'hC60: exp_out = 32'h00174560; // x = -7.2500, f(x) = 0.0007
          12'hC61: exp_out = 32'h00177419; // x = -7.2422, f(x) = 0.0007
          12'hC62: exp_out = 32'h0017A331; // x = -7.2344, f(x) = 0.0007
          12'hC63: exp_out = 32'h0017D2A6; // x = -7.2266, f(x) = 0.0007
          12'hC64: exp_out = 32'h0018027B; // x = -7.2188, f(x) = 0.0007
          12'hC65: exp_out = 32'h001832B0; // x = -7.2109, f(x) = 0.0007
          12'hC66: exp_out = 32'h00186346; // x = -7.2031, f(x) = 0.0007
          12'hC67: exp_out = 32'h0018943E; // x = -7.1953, f(x) = 0.0008
          12'hC68: exp_out = 32'h0018C598; // x = -7.1875, f(x) = 0.0008
          12'hC69: exp_out = 32'h0018F754; // x = -7.1797, f(x) = 0.0008
          12'hC6A: exp_out = 32'h00192975; // x = -7.1719, f(x) = 0.0008
          12'hC6B: exp_out = 32'h00195BFB; // x = -7.1641, f(x) = 0.0008
          12'hC6C: exp_out = 32'h00198EE5; // x = -7.1562, f(x) = 0.0008
          12'hC6D: exp_out = 32'h0019C236; // x = -7.1484, f(x) = 0.0008
          12'hC6E: exp_out = 32'h0019F5EE; // x = -7.1406, f(x) = 0.0008
          12'hC6F: exp_out = 32'h001A2A0E; // x = -7.1328, f(x) = 0.0008
          12'hC70: exp_out = 32'h001A5E97; // x = -7.1250, f(x) = 0.0008
          12'hC71: exp_out = 32'h001A9389; // x = -7.1172, f(x) = 0.0008
          12'hC72: exp_out = 32'h001AC8E5; // x = -7.1094, f(x) = 0.0008
          12'hC73: exp_out = 32'h001AFEAD; // x = -7.1016, f(x) = 0.0008
          12'hC74: exp_out = 32'h001B34E0; // x = -7.0938, f(x) = 0.0008
          12'hC75: exp_out = 32'h001B6B81; // x = -7.0859, f(x) = 0.0008
          12'hC76: exp_out = 32'h001BA28F; // x = -7.0781, f(x) = 0.0008
          12'hC77: exp_out = 32'h001BDA0B; // x = -7.0703, f(x) = 0.0008
          12'hC78: exp_out = 32'h001C11F7; // x = -7.0625, f(x) = 0.0009
          12'hC79: exp_out = 32'h001C4A53; // x = -7.0547, f(x) = 0.0009
          12'hC7A: exp_out = 32'h001C8321; // x = -7.0469, f(x) = 0.0009
          12'hC7B: exp_out = 32'h001CBC60; // x = -7.0391, f(x) = 0.0009
          12'hC7C: exp_out = 32'h001CF613; // x = -7.0312, f(x) = 0.0009
          12'hC7D: exp_out = 32'h001D3039; // x = -7.0234, f(x) = 0.0009
          12'hC7E: exp_out = 32'h001D6AD4; // x = -7.0156, f(x) = 0.0009
          12'hC7F: exp_out = 32'h001DA5E4; // x = -7.0078, f(x) = 0.0009
          12'hC80: exp_out = 32'h001DE16C; // x = -7.0000, f(x) = 0.0009
          12'hC81: exp_out = 32'h001E1D6A; // x = -6.9922, f(x) = 0.0009
          12'hC82: exp_out = 32'h001E59E2; // x = -6.9844, f(x) = 0.0009
          12'hC83: exp_out = 32'h001E96D2; // x = -6.9766, f(x) = 0.0009
          12'hC84: exp_out = 32'h001ED43D; // x = -6.9688, f(x) = 0.0009
          12'hC85: exp_out = 32'h001F1223; // x = -6.9609, f(x) = 0.0009
          12'hC86: exp_out = 32'h001F5086; // x = -6.9531, f(x) = 0.0010
          12'hC87: exp_out = 32'h001F8F66; // x = -6.9453, f(x) = 0.0010
          12'hC88: exp_out = 32'h001FCEC4; // x = -6.9375, f(x) = 0.0010
          12'hC89: exp_out = 32'h00200EA1; // x = -6.9297, f(x) = 0.0010
          12'hC8A: exp_out = 32'h00204EFF; // x = -6.9219, f(x) = 0.0010
          12'hC8B: exp_out = 32'h00208FDE; // x = -6.9141, f(x) = 0.0010
          12'hC8C: exp_out = 32'h0020D13F; // x = -6.9062, f(x) = 0.0010
          12'hC8D: exp_out = 32'h00211323; // x = -6.8984, f(x) = 0.0010
          12'hC8E: exp_out = 32'h0021558C; // x = -6.8906, f(x) = 0.0010
          12'hC8F: exp_out = 32'h00219879; // x = -6.8828, f(x) = 0.0010
          12'hC90: exp_out = 32'h0021DBEE; // x = -6.8750, f(x) = 0.0010
          12'hC91: exp_out = 32'h00221FEA; // x = -6.8672, f(x) = 0.0010
          12'hC92: exp_out = 32'h0022646E; // x = -6.8594, f(x) = 0.0010
          12'hC93: exp_out = 32'h0022A97C; // x = -6.8516, f(x) = 0.0011
          12'hC94: exp_out = 32'h0022EF14; // x = -6.8438, f(x) = 0.0011
          12'hC95: exp_out = 32'h00233538; // x = -6.8359, f(x) = 0.0011
          12'hC96: exp_out = 32'h00237BE9; // x = -6.8281, f(x) = 0.0011
          12'hC97: exp_out = 32'h0023C328; // x = -6.8203, f(x) = 0.0011
          12'hC98: exp_out = 32'h00240AF6; // x = -6.8125, f(x) = 0.0011
          12'hC99: exp_out = 32'h00245355; // x = -6.8047, f(x) = 0.0011
          12'hC9A: exp_out = 32'h00249C44; // x = -6.7969, f(x) = 0.0011
          12'hC9B: exp_out = 32'h0024E5C6; // x = -6.7891, f(x) = 0.0011
          12'hC9C: exp_out = 32'h00252FDC; // x = -6.7812, f(x) = 0.0011
          12'hC9D: exp_out = 32'h00257A86; // x = -6.7734, f(x) = 0.0011
          12'hC9E: exp_out = 32'h0025C5C6; // x = -6.7656, f(x) = 0.0012
          12'hC9F: exp_out = 32'h0026119D; // x = -6.7578, f(x) = 0.0012
          12'hCA0: exp_out = 32'h00265E0D; // x = -6.7500, f(x) = 0.0012
          12'hCA1: exp_out = 32'h0026AB16; // x = -6.7422, f(x) = 0.0012
          12'hCA2: exp_out = 32'h0026F8BA; // x = -6.7344, f(x) = 0.0012
          12'hCA3: exp_out = 32'h002746F9; // x = -6.7266, f(x) = 0.0012
          12'hCA4: exp_out = 32'h002795D6; // x = -6.7188, f(x) = 0.0012
          12'hCA5: exp_out = 32'h0027E551; // x = -6.7109, f(x) = 0.0012
          12'hCA6: exp_out = 32'h0028356C; // x = -6.7031, f(x) = 0.0012
          12'hCA7: exp_out = 32'h00288627; // x = -6.6953, f(x) = 0.0012
          12'hCA8: exp_out = 32'h0028D785; // x = -6.6875, f(x) = 0.0012
          12'hCA9: exp_out = 32'h00292986; // x = -6.6797, f(x) = 0.0013
          12'hCAA: exp_out = 32'h00297C2B; // x = -6.6719, f(x) = 0.0013
          12'hCAB: exp_out = 32'h0029CF77; // x = -6.6641, f(x) = 0.0013
          12'hCAC: exp_out = 32'h002A2369; // x = -6.6562, f(x) = 0.0013
          12'hCAD: exp_out = 32'h002A7805; // x = -6.6484, f(x) = 0.0013
          12'hCAE: exp_out = 32'h002ACD4A; // x = -6.6406, f(x) = 0.0013
          12'hCAF: exp_out = 32'h002B233A; // x = -6.6328, f(x) = 0.0013
          12'hCB0: exp_out = 32'h002B79D7; // x = -6.6250, f(x) = 0.0013
          12'hCB1: exp_out = 32'h002BD122; // x = -6.6172, f(x) = 0.0013
          12'hCB2: exp_out = 32'h002C291C; // x = -6.6094, f(x) = 0.0013
          12'hCB3: exp_out = 32'h002C81C7; // x = -6.6016, f(x) = 0.0014
          12'hCB4: exp_out = 32'h002CDB24; // x = -6.5938, f(x) = 0.0014
          12'hCB5: exp_out = 32'h002D3534; // x = -6.5859, f(x) = 0.0014
          12'hCB6: exp_out = 32'h002D8FF9; // x = -6.5781, f(x) = 0.0014
          12'hCB7: exp_out = 32'h002DEB74; // x = -6.5703, f(x) = 0.0014
          12'hCB8: exp_out = 32'h002E47A7; // x = -6.5625, f(x) = 0.0014
          12'hCB9: exp_out = 32'h002EA494; // x = -6.5547, f(x) = 0.0014
          12'hCBA: exp_out = 32'h002F023A; // x = -6.5469, f(x) = 0.0014
          12'hCBB: exp_out = 32'h002F609D; // x = -6.5391, f(x) = 0.0014
          12'hCBC: exp_out = 32'h002FBFBD; // x = -6.5312, f(x) = 0.0015
          12'hCBD: exp_out = 32'h00301F9C; // x = -6.5234, f(x) = 0.0015
          12'hCBE: exp_out = 32'h0030803C; // x = -6.5156, f(x) = 0.0015
          12'hCBF: exp_out = 32'h0030E19E; // x = -6.5078, f(x) = 0.0015
          12'hCC0: exp_out = 32'h003143C3; // x = -6.5000, f(x) = 0.0015
          12'hCC1: exp_out = 32'h0031A6AD; // x = -6.4922, f(x) = 0.0015
          12'hCC2: exp_out = 32'h00320A5E; // x = -6.4844, f(x) = 0.0015
          12'hCC3: exp_out = 32'h00326ED7; // x = -6.4766, f(x) = 0.0015
          12'hCC4: exp_out = 32'h0032D41A; // x = -6.4688, f(x) = 0.0016
          12'hCC5: exp_out = 32'h00333A28; // x = -6.4609, f(x) = 0.0016
          12'hCC6: exp_out = 32'h0033A103; // x = -6.4531, f(x) = 0.0016
          12'hCC7: exp_out = 32'h003408AD; // x = -6.4453, f(x) = 0.0016
          12'hCC8: exp_out = 32'h00347127; // x = -6.4375, f(x) = 0.0016
          12'hCC9: exp_out = 32'h0034DA72; // x = -6.4297, f(x) = 0.0016
          12'hCCA: exp_out = 32'h00354491; // x = -6.4219, f(x) = 0.0016
          12'hCCB: exp_out = 32'h0035AF85; // x = -6.4141, f(x) = 0.0016
          12'hCCC: exp_out = 32'h00361B50; // x = -6.4062, f(x) = 0.0017
          12'hCCD: exp_out = 32'h003687F3; // x = -6.3984, f(x) = 0.0017
          12'hCCE: exp_out = 32'h0036F570; // x = -6.3906, f(x) = 0.0017
          12'hCCF: exp_out = 32'h003763C9; // x = -6.3828, f(x) = 0.0017
          12'hCD0: exp_out = 32'h0037D300; // x = -6.3750, f(x) = 0.0017
          12'hCD1: exp_out = 32'h00384316; // x = -6.3672, f(x) = 0.0017
          12'hCD2: exp_out = 32'h0038B40D; // x = -6.3594, f(x) = 0.0017
          12'hCD3: exp_out = 32'h003925E6; // x = -6.3516, f(x) = 0.0017
          12'hCD4: exp_out = 32'h003998A5; // x = -6.3438, f(x) = 0.0018
          12'hCD5: exp_out = 32'h003A0C4A; // x = -6.3359, f(x) = 0.0018
          12'hCD6: exp_out = 32'h003A80D7; // x = -6.3281, f(x) = 0.0018
          12'hCD7: exp_out = 32'h003AF64E; // x = -6.3203, f(x) = 0.0018
          12'hCD8: exp_out = 32'h003B6CB0; // x = -6.3125, f(x) = 0.0018
          12'hCD9: exp_out = 32'h003BE401; // x = -6.3047, f(x) = 0.0018
          12'hCDA: exp_out = 32'h003C5C41; // x = -6.2969, f(x) = 0.0018
          12'hCDB: exp_out = 32'h003CD573; // x = -6.2891, f(x) = 0.0019
          12'hCDC: exp_out = 32'h003D4F97; // x = -6.2812, f(x) = 0.0019
          12'hCDD: exp_out = 32'h003DCAB2; // x = -6.2734, f(x) = 0.0019
          12'hCDE: exp_out = 32'h003E46C3; // x = -6.2656, f(x) = 0.0019
          12'hCDF: exp_out = 32'h003EC3CD; // x = -6.2578, f(x) = 0.0019
          12'hCE0: exp_out = 32'h003F41D3; // x = -6.2500, f(x) = 0.0019
          12'hCE1: exp_out = 32'h003FC0D5; // x = -6.2422, f(x) = 0.0019
          12'hCE2: exp_out = 32'h004040D7; // x = -6.2344, f(x) = 0.0020
          12'hCE3: exp_out = 32'h0040C1D9; // x = -6.2266, f(x) = 0.0020
          12'hCE4: exp_out = 32'h004143DF; // x = -6.2188, f(x) = 0.0020
          12'hCE5: exp_out = 32'h0041C6E9; // x = -6.2109, f(x) = 0.0020
          12'hCE6: exp_out = 32'h00424AFB; // x = -6.2031, f(x) = 0.0020
          12'hCE7: exp_out = 32'h0042D016; // x = -6.1953, f(x) = 0.0020
          12'hCE8: exp_out = 32'h0043563C; // x = -6.1875, f(x) = 0.0021
          12'hCE9: exp_out = 32'h0043DD70; // x = -6.1797, f(x) = 0.0021
          12'hCEA: exp_out = 32'h004465B3; // x = -6.1719, f(x) = 0.0021
          12'hCEB: exp_out = 32'h0044EF07; // x = -6.1641, f(x) = 0.0021
          12'hCEC: exp_out = 32'h0045796F; // x = -6.1562, f(x) = 0.0021
          12'hCED: exp_out = 32'h004604EE; // x = -6.1484, f(x) = 0.0021
          12'hCEE: exp_out = 32'h00469184; // x = -6.1406, f(x) = 0.0022
          12'hCEF: exp_out = 32'h00471F34; // x = -6.1328, f(x) = 0.0022
          12'hCF0: exp_out = 32'h0047AE01; // x = -6.1250, f(x) = 0.0022
          12'hCF1: exp_out = 32'h00483DED; // x = -6.1172, f(x) = 0.0022
          12'hCF2: exp_out = 32'h0048CEFA; // x = -6.1094, f(x) = 0.0022
          12'hCF3: exp_out = 32'h0049612A; // x = -6.1016, f(x) = 0.0022
          12'hCF4: exp_out = 32'h0049F47F; // x = -6.0938, f(x) = 0.0023
          12'hCF5: exp_out = 32'h004A88FD; // x = -6.0859, f(x) = 0.0023
          12'hCF6: exp_out = 32'h004B1EA4; // x = -6.0781, f(x) = 0.0023
          12'hCF7: exp_out = 32'h004BB578; // x = -6.0703, f(x) = 0.0023
          12'hCF8: exp_out = 32'h004C4D7B; // x = -6.0625, f(x) = 0.0023
          12'hCF9: exp_out = 32'h004CE6AF; // x = -6.0547, f(x) = 0.0023
          12'hCFA: exp_out = 32'h004D8116; // x = -6.0469, f(x) = 0.0024
          12'hCFB: exp_out = 32'h004E1CB4; // x = -6.0391, f(x) = 0.0024
          12'hCFC: exp_out = 32'h004EB98A; // x = -6.0312, f(x) = 0.0024
          12'hCFD: exp_out = 32'h004F579B; // x = -6.0234, f(x) = 0.0024
          12'hCFE: exp_out = 32'h004FF6E9; // x = -6.0156, f(x) = 0.0024
          12'hCFF: exp_out = 32'h00509777; // x = -6.0078, f(x) = 0.0025
          12'hD00: exp_out = 32'h00513948; // x = -6.0000, f(x) = 0.0025
          12'hD01: exp_out = 32'h0051DC5D; // x = -5.9922, f(x) = 0.0025
          12'hD02: exp_out = 32'h005280BA; // x = -5.9844, f(x) = 0.0025
          12'hD03: exp_out = 32'h00532661; // x = -5.9766, f(x) = 0.0025
          12'hD04: exp_out = 32'h0053CD54; // x = -5.9688, f(x) = 0.0026
          12'hD05: exp_out = 32'h00547597; // x = -5.9609, f(x) = 0.0026
          12'hD06: exp_out = 32'h00551F2C; // x = -5.9531, f(x) = 0.0026
          12'hD07: exp_out = 32'h0055CA15; // x = -5.9453, f(x) = 0.0026
          12'hD08: exp_out = 32'h00567655; // x = -5.9375, f(x) = 0.0026
          12'hD09: exp_out = 32'h005723EF; // x = -5.9297, f(x) = 0.0027
          12'hD0A: exp_out = 32'h0057D2E6; // x = -5.9219, f(x) = 0.0027
          12'hD0B: exp_out = 32'h0058833B; // x = -5.9141, f(x) = 0.0027
          12'hD0C: exp_out = 32'h005934F3; // x = -5.9062, f(x) = 0.0027
          12'hD0D: exp_out = 32'h0059E810; // x = -5.8984, f(x) = 0.0027
          12'hD0E: exp_out = 32'h005A9C95; // x = -5.8906, f(x) = 0.0028
          12'hD0F: exp_out = 32'h005B5283; // x = -5.8828, f(x) = 0.0028
          12'hD10: exp_out = 32'h005C09E0; // x = -5.8750, f(x) = 0.0028
          12'hD11: exp_out = 32'h005CC2AC; // x = -5.8672, f(x) = 0.0028
          12'hD12: exp_out = 32'h005D7CEB; // x = -5.8594, f(x) = 0.0029
          12'hD13: exp_out = 32'h005E38A1; // x = -5.8516, f(x) = 0.0029
          12'hD14: exp_out = 32'h005EF5CF; // x = -5.8438, f(x) = 0.0029
          12'hD15: exp_out = 32'h005FB479; // x = -5.8359, f(x) = 0.0029
          12'hD16: exp_out = 32'h006074A2; // x = -5.8281, f(x) = 0.0029
          12'hD17: exp_out = 32'h0061364C; // x = -5.8203, f(x) = 0.0030
          12'hD18: exp_out = 32'h0061F97C; // x = -5.8125, f(x) = 0.0030
          12'hD19: exp_out = 32'h0062BE33; // x = -5.8047, f(x) = 0.0030
          12'hD1A: exp_out = 32'h00638476; // x = -5.7969, f(x) = 0.0030
          12'hD1B: exp_out = 32'h00644C46; // x = -5.7891, f(x) = 0.0031
          12'hD1C: exp_out = 32'h006515A8; // x = -5.7812, f(x) = 0.0031
          12'hD1D: exp_out = 32'h0065E09E; // x = -5.7734, f(x) = 0.0031
          12'hD1E: exp_out = 32'h0066AD2B; // x = -5.7656, f(x) = 0.0031
          12'hD1F: exp_out = 32'h00677B54; // x = -5.7578, f(x) = 0.0032
          12'hD20: exp_out = 32'h00684B1A; // x = -5.7500, f(x) = 0.0032
          12'hD21: exp_out = 32'h00691C81; // x = -5.7422, f(x) = 0.0032
          12'hD22: exp_out = 32'h0069EF8D; // x = -5.7344, f(x) = 0.0032
          12'hD23: exp_out = 32'h006AC440; // x = -5.7266, f(x) = 0.0033
          12'hD24: exp_out = 32'h006B9A9F; // x = -5.7188, f(x) = 0.0033
          12'hD25: exp_out = 32'h006C72AC; // x = -5.7109, f(x) = 0.0033
          12'hD26: exp_out = 32'h006D4C6B; // x = -5.7031, f(x) = 0.0033
          12'hD27: exp_out = 32'h006E27DF; // x = -5.6953, f(x) = 0.0034
          12'hD28: exp_out = 32'h006F050B; // x = -5.6875, f(x) = 0.0034
          12'hD29: exp_out = 32'h006FE3F4; // x = -5.6797, f(x) = 0.0034
          12'hD2A: exp_out = 32'h0070C49C; // x = -5.6719, f(x) = 0.0034
          12'hD2B: exp_out = 32'h0071A708; // x = -5.6641, f(x) = 0.0035
          12'hD2C: exp_out = 32'h00728B3A; // x = -5.6562, f(x) = 0.0035
          12'hD2D: exp_out = 32'h00737136; // x = -5.6484, f(x) = 0.0035
          12'hD2E: exp_out = 32'h00745900; // x = -5.6406, f(x) = 0.0036
          12'hD2F: exp_out = 32'h0075429B; // x = -5.6328, f(x) = 0.0036
          12'hD30: exp_out = 32'h00762E0B; // x = -5.6250, f(x) = 0.0036
          12'hD31: exp_out = 32'h00771B54; // x = -5.6172, f(x) = 0.0036
          12'hD32: exp_out = 32'h00780A7A; // x = -5.6094, f(x) = 0.0037
          12'hD33: exp_out = 32'h0078FB80; // x = -5.6016, f(x) = 0.0037
          12'hD34: exp_out = 32'h0079EE69; // x = -5.5938, f(x) = 0.0037
          12'hD35: exp_out = 32'h007AE33A; // x = -5.5859, f(x) = 0.0038
          12'hD36: exp_out = 32'h007BD9F7; // x = -5.5781, f(x) = 0.0038
          12'hD37: exp_out = 32'h007CD2A4; // x = -5.5703, f(x) = 0.0038
          12'hD38: exp_out = 32'h007DCD43; // x = -5.5625, f(x) = 0.0038
          12'hD39: exp_out = 32'h007EC9DA; // x = -5.5547, f(x) = 0.0039
          12'hD3A: exp_out = 32'h007FC86C; // x = -5.5469, f(x) = 0.0039
          12'hD3B: exp_out = 32'h0080C8FD; // x = -5.5391, f(x) = 0.0039
          12'hD3C: exp_out = 32'h0081CB91; // x = -5.5312, f(x) = 0.0040
          12'hD3D: exp_out = 32'h0082D02D; // x = -5.5234, f(x) = 0.0040
          12'hD3E: exp_out = 32'h0083D6D3; // x = -5.5156, f(x) = 0.0040
          12'hD3F: exp_out = 32'h0084DF89; // x = -5.5078, f(x) = 0.0041
          12'hD40: exp_out = 32'h0085EA53; // x = -5.5000, f(x) = 0.0041
          12'hD41: exp_out = 32'h0086F734; // x = -5.4922, f(x) = 0.0041
          12'hD42: exp_out = 32'h00880631; // x = -5.4844, f(x) = 0.0042
          12'hD43: exp_out = 32'h0089174E; // x = -5.4766, f(x) = 0.0042
          12'hD44: exp_out = 32'h008A2A90; // x = -5.4688, f(x) = 0.0042
          12'hD45: exp_out = 32'h008B3FFA; // x = -5.4609, f(x) = 0.0042
          12'hD46: exp_out = 32'h008C5791; // x = -5.4531, f(x) = 0.0043
          12'hD47: exp_out = 32'h008D715A; // x = -5.4453, f(x) = 0.0043
          12'hD48: exp_out = 32'h008E8D58; // x = -5.4375, f(x) = 0.0044
          12'hD49: exp_out = 32'h008FAB90; // x = -5.4297, f(x) = 0.0044
          12'hD4A: exp_out = 32'h0090CC08; // x = -5.4219, f(x) = 0.0044
          12'hD4B: exp_out = 32'h0091EEC2; // x = -5.4141, f(x) = 0.0045
          12'hD4C: exp_out = 32'h009313C4; // x = -5.4062, f(x) = 0.0045
          12'hD4D: exp_out = 32'h00943B13; // x = -5.3984, f(x) = 0.0045
          12'hD4E: exp_out = 32'h009564B2; // x = -5.3906, f(x) = 0.0046
          12'hD4F: exp_out = 32'h009690A7; // x = -5.3828, f(x) = 0.0046
          12'hD50: exp_out = 32'h0097BEF6; // x = -5.3750, f(x) = 0.0046
          12'hD51: exp_out = 32'h0098EFA4; // x = -5.3672, f(x) = 0.0047
          12'hD52: exp_out = 32'h009A22B6; // x = -5.3594, f(x) = 0.0047
          12'hD53: exp_out = 32'h009B5831; // x = -5.3516, f(x) = 0.0047
          12'hD54: exp_out = 32'h009C9019; // x = -5.3438, f(x) = 0.0048
          12'hD55: exp_out = 32'h009DCA73; // x = -5.3359, f(x) = 0.0048
          12'hD56: exp_out = 32'h009F0744; // x = -5.3281, f(x) = 0.0049
          12'hD57: exp_out = 32'h00A04692; // x = -5.3203, f(x) = 0.0049
          12'hD58: exp_out = 32'h00A18860; // x = -5.3125, f(x) = 0.0049
          12'hD59: exp_out = 32'h00A2CCB5; // x = -5.3047, f(x) = 0.0050
          12'hD5A: exp_out = 32'h00A41395; // x = -5.2969, f(x) = 0.0050
          12'hD5B: exp_out = 32'h00A55D05; // x = -5.2891, f(x) = 0.0050
          12'hD5C: exp_out = 32'h00A6A90B; // x = -5.2812, f(x) = 0.0051
          12'hD5D: exp_out = 32'h00A7F7AB; // x = -5.2734, f(x) = 0.0051
          12'hD5E: exp_out = 32'h00A948EB; // x = -5.2656, f(x) = 0.0052
          12'hD5F: exp_out = 32'h00AA9CD0; // x = -5.2578, f(x) = 0.0052
          12'hD60: exp_out = 32'h00ABF360; // x = -5.2500, f(x) = 0.0052
          12'hD61: exp_out = 32'h00AD4CA0; // x = -5.2422, f(x) = 0.0053
          12'hD62: exp_out = 32'h00AEA894; // x = -5.2344, f(x) = 0.0053
          12'hD63: exp_out = 32'h00B00744; // x = -5.2266, f(x) = 0.0054
          12'hD64: exp_out = 32'h00B168B3; // x = -5.2188, f(x) = 0.0054
          12'hD65: exp_out = 32'h00B2CCE8; // x = -5.2109, f(x) = 0.0055
          12'hD66: exp_out = 32'h00B433E9; // x = -5.2031, f(x) = 0.0055
          12'hD67: exp_out = 32'h00B59DBA; // x = -5.1953, f(x) = 0.0055
          12'hD68: exp_out = 32'h00B70A61; // x = -5.1875, f(x) = 0.0056
          12'hD69: exp_out = 32'h00B879E5; // x = -5.1797, f(x) = 0.0056
          12'hD6A: exp_out = 32'h00B9EC4B; // x = -5.1719, f(x) = 0.0057
          12'hD6B: exp_out = 32'h00BB6198; // x = -5.1641, f(x) = 0.0057
          12'hD6C: exp_out = 32'h00BCD9D3; // x = -5.1562, f(x) = 0.0058
          12'hD6D: exp_out = 32'h00BE5502; // x = -5.1484, f(x) = 0.0058
          12'hD6E: exp_out = 32'h00BFD329; // x = -5.1406, f(x) = 0.0059
          12'hD6F: exp_out = 32'h00C15450; // x = -5.1328, f(x) = 0.0059
          12'hD70: exp_out = 32'h00C2D87D; // x = -5.1250, f(x) = 0.0059
          12'hD71: exp_out = 32'h00C45FB4; // x = -5.1172, f(x) = 0.0060
          12'hD72: exp_out = 32'h00C5E9FD; // x = -5.1094, f(x) = 0.0060
          12'hD73: exp_out = 32'h00C7775E; // x = -5.1016, f(x) = 0.0061
          12'hD74: exp_out = 32'h00C907DD; // x = -5.0938, f(x) = 0.0061
          12'hD75: exp_out = 32'h00CA9B80; // x = -5.0859, f(x) = 0.0062
          12'hD76: exp_out = 32'h00CC324D; // x = -5.0781, f(x) = 0.0062
          12'hD77: exp_out = 32'h00CDCC4B; // x = -5.0703, f(x) = 0.0063
          12'hD78: exp_out = 32'h00CF6980; // x = -5.0625, f(x) = 0.0063
          12'hD79: exp_out = 32'h00D109F3; // x = -5.0547, f(x) = 0.0064
          12'hD7A: exp_out = 32'h00D2ADAA; // x = -5.0469, f(x) = 0.0064
          12'hD7B: exp_out = 32'h00D454AC; // x = -5.0391, f(x) = 0.0065
          12'hD7C: exp_out = 32'h00D5FEFF; // x = -5.0312, f(x) = 0.0065
          12'hD7D: exp_out = 32'h00D7ACAA; // x = -5.0234, f(x) = 0.0066
          12'hD7E: exp_out = 32'h00D95DB4; // x = -5.0156, f(x) = 0.0066
          12'hD7F: exp_out = 32'h00DB1223; // x = -5.0078, f(x) = 0.0067
          12'hD80: exp_out = 32'h00DCC9FF; // x = -5.0000, f(x) = 0.0067
          12'hD81: exp_out = 32'h00DE854E; // x = -4.9922, f(x) = 0.0068
          12'hD82: exp_out = 32'h00E04417; // x = -4.9844, f(x) = 0.0068
          12'hD83: exp_out = 32'h00E20660; // x = -4.9766, f(x) = 0.0069
          12'hD84: exp_out = 32'h00E3CC32; // x = -4.9688, f(x) = 0.0070
          12'hD85: exp_out = 32'h00E59594; // x = -4.9609, f(x) = 0.0070
          12'hD86: exp_out = 32'h00E7628B; // x = -4.9531, f(x) = 0.0071
          12'hD87: exp_out = 32'h00E93320; // x = -4.9453, f(x) = 0.0071
          12'hD88: exp_out = 32'h00EB075A; // x = -4.9375, f(x) = 0.0072
          12'hD89: exp_out = 32'h00ECDF40; // x = -4.9297, f(x) = 0.0072
          12'hD8A: exp_out = 32'h00EEBAD9; // x = -4.9219, f(x) = 0.0073
          12'hD8B: exp_out = 32'h00F09A2E; // x = -4.9141, f(x) = 0.0073
          12'hD8C: exp_out = 32'h00F27D45; // x = -4.9062, f(x) = 0.0074
          12'hD8D: exp_out = 32'h00F46425; // x = -4.8984, f(x) = 0.0075
          12'hD8E: exp_out = 32'h00F64ED8; // x = -4.8906, f(x) = 0.0075
          12'hD8F: exp_out = 32'h00F83D63; // x = -4.8828, f(x) = 0.0076
          12'hD90: exp_out = 32'h00FA2FD0; // x = -4.8750, f(x) = 0.0076
          12'hD91: exp_out = 32'h00FC2625; // x = -4.8672, f(x) = 0.0077
          12'hD92: exp_out = 32'h00FE206B; // x = -4.8594, f(x) = 0.0078
          12'hD93: exp_out = 32'h01001EAA; // x = -4.8516, f(x) = 0.0078
          12'hD94: exp_out = 32'h010220E9; // x = -4.8438, f(x) = 0.0079
          12'hD95: exp_out = 32'h01042730; // x = -4.8359, f(x) = 0.0079
          12'hD96: exp_out = 32'h01063188; // x = -4.8281, f(x) = 0.0080
          12'hD97: exp_out = 32'h01083FF9; // x = -4.8203, f(x) = 0.0081
          12'hD98: exp_out = 32'h010A528B; // x = -4.8125, f(x) = 0.0081
          12'hD99: exp_out = 32'h010C6946; // x = -4.8047, f(x) = 0.0082
          12'hD9A: exp_out = 32'h010E8432; // x = -4.7969, f(x) = 0.0083
          12'hD9B: exp_out = 32'h0110A359; // x = -4.7891, f(x) = 0.0083
          12'hD9C: exp_out = 32'h0112C6C3; // x = -4.7812, f(x) = 0.0084
          12'hD9D: exp_out = 32'h0114EE77; // x = -4.7734, f(x) = 0.0085
          12'hD9E: exp_out = 32'h01171A7F; // x = -4.7656, f(x) = 0.0085
          12'hD9F: exp_out = 32'h01194AE4; // x = -4.7578, f(x) = 0.0086
          12'hDA0: exp_out = 32'h011B7FAE; // x = -4.7500, f(x) = 0.0087
          12'hDA1: exp_out = 32'h011DB8E6; // x = -4.7422, f(x) = 0.0087
          12'hDA2: exp_out = 32'h011FF695; // x = -4.7344, f(x) = 0.0088
          12'hDA3: exp_out = 32'h012238C3; // x = -4.7266, f(x) = 0.0089
          12'hDA4: exp_out = 32'h01247F7B; // x = -4.7188, f(x) = 0.0089
          12'hDA5: exp_out = 32'h0126CAC4; // x = -4.7109, f(x) = 0.0090
          12'hDA6: exp_out = 32'h01291AA9; // x = -4.7031, f(x) = 0.0091
          12'hDA7: exp_out = 32'h012B6F32; // x = -4.6953, f(x) = 0.0091
          12'hDA8: exp_out = 32'h012DC869; // x = -4.6875, f(x) = 0.0092
          12'hDA9: exp_out = 32'h01302657; // x = -4.6797, f(x) = 0.0093
          12'hDAA: exp_out = 32'h01328905; // x = -4.6719, f(x) = 0.0094
          12'hDAB: exp_out = 32'h0134F07E; // x = -4.6641, f(x) = 0.0094
          12'hDAC: exp_out = 32'h01375CCA; // x = -4.6562, f(x) = 0.0095
          12'hDAD: exp_out = 32'h0139CDF4; // x = -4.6484, f(x) = 0.0096
          12'hDAE: exp_out = 32'h013C4405; // x = -4.6406, f(x) = 0.0097
          12'hDAF: exp_out = 32'h013EBF08; // x = -4.6328, f(x) = 0.0097
          12'hDB0: exp_out = 32'h01413F05; // x = -4.6250, f(x) = 0.0098
          12'hDB1: exp_out = 32'h0143C407; // x = -4.6172, f(x) = 0.0099
          12'hDB2: exp_out = 32'h01464E18; // x = -4.6094, f(x) = 0.0100
          12'hDB3: exp_out = 32'h0148DD43; // x = -4.6016, f(x) = 0.0100
          12'hDB4: exp_out = 32'h014B7191; // x = -4.5938, f(x) = 0.0101
          12'hDB5: exp_out = 32'h014E0B0D; // x = -4.5859, f(x) = 0.0102
          12'hDB6: exp_out = 32'h0150A9C1; // x = -4.5781, f(x) = 0.0103
          12'hDB7: exp_out = 32'h01534DB7; // x = -4.5703, f(x) = 0.0104
          12'hDB8: exp_out = 32'h0155F6FB; // x = -4.5625, f(x) = 0.0104
          12'hDB9: exp_out = 32'h0158A597; // x = -4.5547, f(x) = 0.0105
          12'hDBA: exp_out = 32'h015B5995; // x = -4.5469, f(x) = 0.0106
          12'hDBB: exp_out = 32'h015E1301; // x = -4.5391, f(x) = 0.0107
          12'hDBC: exp_out = 32'h0160D1E5; // x = -4.5312, f(x) = 0.0108
          12'hDBD: exp_out = 32'h0163964C; // x = -4.5234, f(x) = 0.0109
          12'hDBE: exp_out = 32'h01666041; // x = -4.5156, f(x) = 0.0109
          12'hDBF: exp_out = 32'h01692FD1; // x = -4.5078, f(x) = 0.0110
          12'hDC0: exp_out = 32'h016C0504; // x = -4.5000, f(x) = 0.0111
          12'hDC1: exp_out = 32'h016EDFE8; // x = -4.4922, f(x) = 0.0112
          12'hDC2: exp_out = 32'h0171C088; // x = -4.4844, f(x) = 0.0113
          12'hDC3: exp_out = 32'h0174A6EE; // x = -4.4766, f(x) = 0.0114
          12'hDC4: exp_out = 32'h01779327; // x = -4.4688, f(x) = 0.0115
          12'hDC5: exp_out = 32'h017A853F; // x = -4.4609, f(x) = 0.0116
          12'hDC6: exp_out = 32'h017D7D40; // x = -4.4531, f(x) = 0.0116
          12'hDC7: exp_out = 32'h01807B38; // x = -4.4453, f(x) = 0.0117
          12'hDC8: exp_out = 32'h01837F31; // x = -4.4375, f(x) = 0.0118
          12'hDC9: exp_out = 32'h01868939; // x = -4.4297, f(x) = 0.0119
          12'hDCA: exp_out = 32'h0189995A; // x = -4.4219, f(x) = 0.0120
          12'hDCB: exp_out = 32'h018CAFA2; // x = -4.4141, f(x) = 0.0121
          12'hDCC: exp_out = 32'h018FCC1D; // x = -4.4062, f(x) = 0.0122
          12'hDCD: exp_out = 32'h0192EED7; // x = -4.3984, f(x) = 0.0123
          12'hDCE: exp_out = 32'h019617DC; // x = -4.3906, f(x) = 0.0124
          12'hDCF: exp_out = 32'h0199473A; // x = -4.3828, f(x) = 0.0125
          12'hDD0: exp_out = 32'h019C7CFE; // x = -4.3750, f(x) = 0.0126
          12'hDD1: exp_out = 32'h019FB933; // x = -4.3672, f(x) = 0.0127
          12'hDD2: exp_out = 32'h01A2FBE7; // x = -4.3594, f(x) = 0.0128
          12'hDD3: exp_out = 32'h01A64527; // x = -4.3516, f(x) = 0.0129
          12'hDD4: exp_out = 32'h01A99500; // x = -4.3438, f(x) = 0.0130
          12'hDD5: exp_out = 32'h01ACEB7F; // x = -4.3359, f(x) = 0.0131
          12'hDD6: exp_out = 32'h01B048B2; // x = -4.3281, f(x) = 0.0132
          12'hDD7: exp_out = 32'h01B3ACA6; // x = -4.3203, f(x) = 0.0133
          12'hDD8: exp_out = 32'h01B71769; // x = -4.3125, f(x) = 0.0134
          12'hDD9: exp_out = 32'h01BA8909; // x = -4.3047, f(x) = 0.0135
          12'hDDA: exp_out = 32'h01BE0192; // x = -4.2969, f(x) = 0.0136
          12'hDDB: exp_out = 32'h01C18114; // x = -4.2891, f(x) = 0.0137
          12'hDDC: exp_out = 32'h01C5079B; // x = -4.2812, f(x) = 0.0138
          12'hDDD: exp_out = 32'h01C89537; // x = -4.2734, f(x) = 0.0139
          12'hDDE: exp_out = 32'h01CC29F5; // x = -4.2656, f(x) = 0.0140
          12'hDDF: exp_out = 32'h01CFC5E3; // x = -4.2578, f(x) = 0.0142
          12'hDE0: exp_out = 32'h01D36911; // x = -4.2500, f(x) = 0.0143
          12'hDE1: exp_out = 32'h01D7138C; // x = -4.2422, f(x) = 0.0144
          12'hDE2: exp_out = 32'h01DAC564; // x = -4.2344, f(x) = 0.0145
          12'hDE3: exp_out = 32'h01DE7EA7; // x = -4.2266, f(x) = 0.0146
          12'hDE4: exp_out = 32'h01E23F64; // x = -4.2188, f(x) = 0.0147
          12'hDE5: exp_out = 32'h01E607AA; // x = -4.2109, f(x) = 0.0148
          12'hDE6: exp_out = 32'h01E9D787; // x = -4.2031, f(x) = 0.0149
          12'hDE7: exp_out = 32'h01EDAF0D; // x = -4.1953, f(x) = 0.0151
          12'hDE8: exp_out = 32'h01F18E49; // x = -4.1875, f(x) = 0.0152
          12'hDE9: exp_out = 32'h01F5754B; // x = -4.1797, f(x) = 0.0153
          12'hDEA: exp_out = 32'h01F96423; // x = -4.1719, f(x) = 0.0154
          12'hDEB: exp_out = 32'h01FD5AE1; // x = -4.1641, f(x) = 0.0155
          12'hDEC: exp_out = 32'h02015994; // x = -4.1562, f(x) = 0.0157
          12'hDED: exp_out = 32'h0205604D; // x = -4.1484, f(x) = 0.0158
          12'hDEE: exp_out = 32'h02096F1B; // x = -4.1406, f(x) = 0.0159
          12'hDEF: exp_out = 32'h020D860E; // x = -4.1328, f(x) = 0.0160
          12'hDF0: exp_out = 32'h0211A538; // x = -4.1250, f(x) = 0.0162
          12'hDF1: exp_out = 32'h0215CCA9; // x = -4.1172, f(x) = 0.0163
          12'hDF2: exp_out = 32'h0219FC71; // x = -4.1094, f(x) = 0.0164
          12'hDF3: exp_out = 32'h021E34A0; // x = -4.1016, f(x) = 0.0165
          12'hDF4: exp_out = 32'h02227549; // x = -4.0938, f(x) = 0.0167
          12'hDF5: exp_out = 32'h0226BE7B; // x = -4.0859, f(x) = 0.0168
          12'hDF6: exp_out = 32'h022B1048; // x = -4.0781, f(x) = 0.0169
          12'hDF7: exp_out = 32'h022F6AC2; // x = -4.0703, f(x) = 0.0171
          12'hDF8: exp_out = 32'h0233CDF9; // x = -4.0625, f(x) = 0.0172
          12'hDF9: exp_out = 32'h02383A00; // x = -4.0547, f(x) = 0.0173
          12'hDFA: exp_out = 32'h023CAEE7; // x = -4.0469, f(x) = 0.0175
          12'hDFB: exp_out = 32'h02412CC1; // x = -4.0391, f(x) = 0.0176
          12'hDFC: exp_out = 32'h0245B3A0; // x = -4.0312, f(x) = 0.0178
          12'hDFD: exp_out = 32'h024A4396; // x = -4.0234, f(x) = 0.0179
          12'hDFE: exp_out = 32'h024EDCB5; // x = -4.0156, f(x) = 0.0180
          12'hDFF: exp_out = 32'h02537F0F; // x = -4.0078, f(x) = 0.0182
          12'hE00: exp_out = 32'h02582AB7; // x = -4.0000, f(x) = 0.0183
          12'hE01: exp_out = 32'h025CDFC0; // x = -3.9922, f(x) = 0.0185
          12'hE02: exp_out = 32'h02619E3C; // x = -3.9844, f(x) = 0.0186
          12'hE03: exp_out = 32'h0266663F; // x = -3.9766, f(x) = 0.0187
          12'hE04: exp_out = 32'h026B37DC; // x = -3.9688, f(x) = 0.0189
          12'hE05: exp_out = 32'h02701325; // x = -3.9609, f(x) = 0.0190
          12'hE06: exp_out = 32'h0274F82F; // x = -3.9531, f(x) = 0.0192
          12'hE07: exp_out = 32'h0279E70C; // x = -3.9453, f(x) = 0.0193
          12'hE08: exp_out = 32'h027EDFD2; // x = -3.9375, f(x) = 0.0195
          12'hE09: exp_out = 32'h0283E292; // x = -3.9297, f(x) = 0.0196
          12'hE0A: exp_out = 32'h0288EF63; // x = -3.9219, f(x) = 0.0198
          12'hE0B: exp_out = 32'h028E0657; // x = -3.9141, f(x) = 0.0200
          12'hE0C: exp_out = 32'h02932783; // x = -3.9062, f(x) = 0.0201
          12'hE0D: exp_out = 32'h029852FC; // x = -3.8984, f(x) = 0.0203
          12'hE0E: exp_out = 32'h029D88D6; // x = -3.8906, f(x) = 0.0204
          12'hE0F: exp_out = 32'h02A2C926; // x = -3.8828, f(x) = 0.0206
          12'hE10: exp_out = 32'h02A81401; // x = -3.8750, f(x) = 0.0208
          12'hE11: exp_out = 32'h02AD697D; // x = -3.8672, f(x) = 0.0209
          12'hE12: exp_out = 32'h02B2C9AE; // x = -3.8594, f(x) = 0.0211
          12'hE13: exp_out = 32'h02B834AB; // x = -3.8516, f(x) = 0.0212
          12'hE14: exp_out = 32'h02BDAA88; // x = -3.8438, f(x) = 0.0214
          12'hE15: exp_out = 32'h02C32B5C; // x = -3.8359, f(x) = 0.0216
          12'hE16: exp_out = 32'h02C8B73D; // x = -3.8281, f(x) = 0.0218
          12'hE17: exp_out = 32'h02CE4E41; // x = -3.8203, f(x) = 0.0219
          12'hE18: exp_out = 32'h02D3F07E; // x = -3.8125, f(x) = 0.0221
          12'hE19: exp_out = 32'h02D99E0A; // x = -3.8047, f(x) = 0.0223
          12'hE1A: exp_out = 32'h02DF56FD; // x = -3.7969, f(x) = 0.0224
          12'hE1B: exp_out = 32'h02E51B6E; // x = -3.7891, f(x) = 0.0226
          12'hE1C: exp_out = 32'h02EAEB73; // x = -3.7812, f(x) = 0.0228
          12'hE1D: exp_out = 32'h02F0C723; // x = -3.7734, f(x) = 0.0230
          12'hE1E: exp_out = 32'h02F6AE97; // x = -3.7656, f(x) = 0.0232
          12'hE1F: exp_out = 32'h02FCA1E6; // x = -3.7578, f(x) = 0.0233
          12'hE20: exp_out = 32'h0302A127; // x = -3.7500, f(x) = 0.0235
          12'hE21: exp_out = 32'h0308AC72; // x = -3.7422, f(x) = 0.0237
          12'hE22: exp_out = 32'h030EC3E1; // x = -3.7344, f(x) = 0.0239
          12'hE23: exp_out = 32'h0314E78A; // x = -3.7266, f(x) = 0.0241
          12'hE24: exp_out = 32'h031B1787; // x = -3.7188, f(x) = 0.0243
          12'hE25: exp_out = 32'h032153F0; // x = -3.7109, f(x) = 0.0245
          12'hE26: exp_out = 32'h03279CDF; // x = -3.7031, f(x) = 0.0246
          12'hE27: exp_out = 32'h032DF26C; // x = -3.6953, f(x) = 0.0248
          12'hE28: exp_out = 32'h033454B1; // x = -3.6875, f(x) = 0.0250
          12'hE29: exp_out = 32'h033AC3C8; // x = -3.6797, f(x) = 0.0252
          12'hE2A: exp_out = 32'h03413FC9; // x = -3.6719, f(x) = 0.0254
          12'hE2B: exp_out = 32'h0347C8CF; // x = -3.6641, f(x) = 0.0256
          12'hE2C: exp_out = 32'h034E5EF5; // x = -3.6562, f(x) = 0.0258
          12'hE2D: exp_out = 32'h03550254; // x = -3.6484, f(x) = 0.0260
          12'hE2E: exp_out = 32'h035BB307; // x = -3.6406, f(x) = 0.0262
          12'hE2F: exp_out = 32'h03627129; // x = -3.6328, f(x) = 0.0264
          12'hE30: exp_out = 32'h03693CD5; // x = -3.6250, f(x) = 0.0266
          12'hE31: exp_out = 32'h03701625; // x = -3.6172, f(x) = 0.0269
          12'hE32: exp_out = 32'h0376FD37; // x = -3.6094, f(x) = 0.0271
          12'hE33: exp_out = 32'h037DF224; // x = -3.6016, f(x) = 0.0273
          12'hE34: exp_out = 32'h0384F508; // x = -3.5938, f(x) = 0.0275
          12'hE35: exp_out = 32'h038C0601; // x = -3.5859, f(x) = 0.0277
          12'hE36: exp_out = 32'h0393252A; // x = -3.5781, f(x) = 0.0279
          12'hE37: exp_out = 32'h039A529F; // x = -3.5703, f(x) = 0.0281
          12'hE38: exp_out = 32'h03A18E7E; // x = -3.5625, f(x) = 0.0284
          12'hE39: exp_out = 32'h03A8D8E3; // x = -3.5547, f(x) = 0.0286
          12'hE3A: exp_out = 32'h03B031EB; // x = -3.5469, f(x) = 0.0288
          12'hE3B: exp_out = 32'h03B799B4; // x = -3.5391, f(x) = 0.0290
          12'hE3C: exp_out = 32'h03BF105C; // x = -3.5312, f(x) = 0.0293
          12'hE3D: exp_out = 32'h03C69600; // x = -3.5234, f(x) = 0.0295
          12'hE3E: exp_out = 32'h03CE2ABE; // x = -3.5156, f(x) = 0.0297
          12'hE3F: exp_out = 32'h03D5CEB5; // x = -3.5078, f(x) = 0.0300
          12'hE40: exp_out = 32'h03DD8203; // x = -3.5000, f(x) = 0.0302
          12'hE41: exp_out = 32'h03E544C7; // x = -3.4922, f(x) = 0.0304
          12'hE42: exp_out = 32'h03ED1721; // x = -3.4844, f(x) = 0.0307
          12'hE43: exp_out = 32'h03F4F92E; // x = -3.4766, f(x) = 0.0309
          12'hE44: exp_out = 32'h03FCEB10; // x = -3.4688, f(x) = 0.0312
          12'hE45: exp_out = 32'h0404ECE5; // x = -3.4609, f(x) = 0.0314
          12'hE46: exp_out = 32'h040CFECE; // x = -3.4531, f(x) = 0.0316
          12'hE47: exp_out = 32'h041520EB; // x = -3.4453, f(x) = 0.0319
          12'hE48: exp_out = 32'h041D535D; // x = -3.4375, f(x) = 0.0321
          12'hE49: exp_out = 32'h04259644; // x = -3.4297, f(x) = 0.0324
          12'hE4A: exp_out = 32'h042DE9C1; // x = -3.4219, f(x) = 0.0327
          12'hE4B: exp_out = 32'h04364DF6; // x = -3.4141, f(x) = 0.0329
          12'hE4C: exp_out = 32'h043EC304; // x = -3.4062, f(x) = 0.0332
          12'hE4D: exp_out = 32'h0447490D; // x = -3.3984, f(x) = 0.0334
          12'hE4E: exp_out = 32'h044FE034; // x = -3.3906, f(x) = 0.0337
          12'hE4F: exp_out = 32'h04588899; // x = -3.3828, f(x) = 0.0340
          12'hE50: exp_out = 32'h04614262; // x = -3.3750, f(x) = 0.0342
          12'hE51: exp_out = 32'h046A0DAF; // x = -3.3672, f(x) = 0.0345
          12'hE52: exp_out = 32'h0472EAA4; // x = -3.3594, f(x) = 0.0348
          12'hE53: exp_out = 32'h047BD965; // x = -3.3516, f(x) = 0.0350
          12'hE54: exp_out = 32'h0484DA16; // x = -3.3438, f(x) = 0.0353
          12'hE55: exp_out = 32'h048DECD9; // x = -3.3359, f(x) = 0.0356
          12'hE56: exp_out = 32'h049711D5; // x = -3.3281, f(x) = 0.0359
          12'hE57: exp_out = 32'h04A0492D; // x = -3.3203, f(x) = 0.0361
          12'hE58: exp_out = 32'h04A99306; // x = -3.3125, f(x) = 0.0364
          12'hE59: exp_out = 32'h04B2EF86; // x = -3.3047, f(x) = 0.0367
          12'hE5A: exp_out = 32'h04BC5ED1; // x = -3.2969, f(x) = 0.0370
          12'hE5B: exp_out = 32'h04C5E10D; // x = -3.2891, f(x) = 0.0373
          12'hE5C: exp_out = 32'h04CF7662; // x = -3.2812, f(x) = 0.0376
          12'hE5D: exp_out = 32'h04D91EF4; // x = -3.2734, f(x) = 0.0379
          12'hE5E: exp_out = 32'h04E2DAEA; // x = -3.2656, f(x) = 0.0382
          12'hE5F: exp_out = 32'h04ECAA6D; // x = -3.2578, f(x) = 0.0385
          12'hE60: exp_out = 32'h04F68DA1; // x = -3.2500, f(x) = 0.0388
          12'hE61: exp_out = 32'h050084B0; // x = -3.2422, f(x) = 0.0391
          12'hE62: exp_out = 32'h050A8FC1; // x = -3.2344, f(x) = 0.0394
          12'hE63: exp_out = 32'h0514AEFD; // x = -3.2266, f(x) = 0.0397
          12'hE64: exp_out = 32'h051EE28B; // x = -3.2188, f(x) = 0.0400
          12'hE65: exp_out = 32'h05292A95; // x = -3.2109, f(x) = 0.0403
          12'hE66: exp_out = 32'h05338743; // x = -3.2031, f(x) = 0.0406
          12'hE67: exp_out = 32'h053DF8BF; // x = -3.1953, f(x) = 0.0410
          12'hE68: exp_out = 32'h05487F34; // x = -3.1875, f(x) = 0.0413
          12'hE69: exp_out = 32'h05531ACA; // x = -3.1797, f(x) = 0.0416
          12'hE6A: exp_out = 32'h055DCBAD; // x = -3.1719, f(x) = 0.0419
          12'hE6B: exp_out = 32'h05689207; // x = -3.1641, f(x) = 0.0423
          12'hE6C: exp_out = 32'h05736E04; // x = -3.1562, f(x) = 0.0426
          12'hE6D: exp_out = 32'h057E5FCE; // x = -3.1484, f(x) = 0.0429
          12'hE6E: exp_out = 32'h05896792; // x = -3.1406, f(x) = 0.0433
          12'hE6F: exp_out = 32'h0594857B; // x = -3.1328, f(x) = 0.0436
          12'hE70: exp_out = 32'h059FB9B6; // x = -3.1250, f(x) = 0.0439
          12'hE71: exp_out = 32'h05AB0471; // x = -3.1172, f(x) = 0.0443
          12'hE72: exp_out = 32'h05B665D7; // x = -3.1094, f(x) = 0.0446
          12'hE73: exp_out = 32'h05C1DE17; // x = -3.1016, f(x) = 0.0450
          12'hE74: exp_out = 32'h05CD6D5F; // x = -3.0938, f(x) = 0.0453
          12'hE75: exp_out = 32'h05D913DC; // x = -3.0859, f(x) = 0.0457
          12'hE76: exp_out = 32'h05E4D1BE; // x = -3.0781, f(x) = 0.0460
          12'hE77: exp_out = 32'h05F0A733; // x = -3.0703, f(x) = 0.0464
          12'hE78: exp_out = 32'h05FC946B; // x = -3.0625, f(x) = 0.0468
          12'hE79: exp_out = 32'h06089995; // x = -3.0547, f(x) = 0.0471
          12'hE7A: exp_out = 32'h0614B6E1; // x = -3.0469, f(x) = 0.0475
          12'hE7B: exp_out = 32'h0620EC81; // x = -3.0391, f(x) = 0.0479
          12'hE7C: exp_out = 32'h062D3AA4; // x = -3.0312, f(x) = 0.0483
          12'hE7D: exp_out = 32'h0639A17C; // x = -3.0234, f(x) = 0.0486
          12'hE7E: exp_out = 32'h0646213A; // x = -3.0156, f(x) = 0.0490
          12'hE7F: exp_out = 32'h0652BA11; // x = -3.0078, f(x) = 0.0494
          12'hE80: exp_out = 32'h065F6C33; // x = -3.0000, f(x) = 0.0498
          12'hE81: exp_out = 32'h066C37D3; // x = -2.9922, f(x) = 0.0502
          12'hE82: exp_out = 32'h06791D24; // x = -2.9844, f(x) = 0.0506
          12'hE83: exp_out = 32'h06861C59; // x = -2.9766, f(x) = 0.0510
          12'hE84: exp_out = 32'h069335A6; // x = -2.9688, f(x) = 0.0514
          12'hE85: exp_out = 32'h06A06941; // x = -2.9609, f(x) = 0.0518
          12'hE86: exp_out = 32'h06ADB75D; // x = -2.9531, f(x) = 0.0522
          12'hE87: exp_out = 32'h06BB2030; // x = -2.9453, f(x) = 0.0526
          12'hE88: exp_out = 32'h06C8A3F0; // x = -2.9375, f(x) = 0.0530
          12'hE89: exp_out = 32'h06D642D2; // x = -2.9297, f(x) = 0.0534
          12'hE8A: exp_out = 32'h06E3FD0D; // x = -2.9219, f(x) = 0.0538
          12'hE8B: exp_out = 32'h06F1D2D9; // x = -2.9141, f(x) = 0.0543
          12'hE8C: exp_out = 32'h06FFC46B; // x = -2.9062, f(x) = 0.0547
          12'hE8D: exp_out = 32'h070DD1FD; // x = -2.8984, f(x) = 0.0551
          12'hE8E: exp_out = 32'h071BFBC6; // x = -2.8906, f(x) = 0.0555
          12'hE8F: exp_out = 32'h072A41FF; // x = -2.8828, f(x) = 0.0560
          12'hE90: exp_out = 32'h0738A4E1; // x = -2.8750, f(x) = 0.0564
          12'hE91: exp_out = 32'h074724A6; // x = -2.8672, f(x) = 0.0569
          12'hE92: exp_out = 32'h0755C187; // x = -2.8594, f(x) = 0.0573
          12'hE93: exp_out = 32'h07647BBF; // x = -2.8516, f(x) = 0.0578
          12'hE94: exp_out = 32'h0773538A; // x = -2.8438, f(x) = 0.0582
          12'hE95: exp_out = 32'h07824921; // x = -2.8359, f(x) = 0.0587
          12'hE96: exp_out = 32'h07915CC2; // x = -2.8281, f(x) = 0.0591
          12'hE97: exp_out = 32'h07A08EA9; // x = -2.8203, f(x) = 0.0596
          12'hE98: exp_out = 32'h07AFDF11; // x = -2.8125, f(x) = 0.0601
          12'hE99: exp_out = 32'h07BF4E39; // x = -2.8047, f(x) = 0.0605
          12'hE9A: exp_out = 32'h07CEDC5F; // x = -2.7969, f(x) = 0.0610
          12'hE9B: exp_out = 32'h07DE89C0; // x = -2.7891, f(x) = 0.0615
          12'hE9C: exp_out = 32'h07EE569B; // x = -2.7812, f(x) = 0.0620
          12'hE9D: exp_out = 32'h07FE432F; // x = -2.7734, f(x) = 0.0624
          12'hE9E: exp_out = 32'h080E4FBD; // x = -2.7656, f(x) = 0.0629
          12'hE9F: exp_out = 32'h081E7C84; // x = -2.7578, f(x) = 0.0634
          12'hEA0: exp_out = 32'h082EC9C5; // x = -2.7500, f(x) = 0.0639
          12'hEA1: exp_out = 32'h083F37C1; // x = -2.7422, f(x) = 0.0644
          12'hEA2: exp_out = 32'h084FC6BA; // x = -2.7344, f(x) = 0.0649
          12'hEA3: exp_out = 32'h086076F2; // x = -2.7266, f(x) = 0.0654
          12'hEA4: exp_out = 32'h087148AC; // x = -2.7188, f(x) = 0.0660
          12'hEA5: exp_out = 32'h08823C2B; // x = -2.7109, f(x) = 0.0665
          12'hEA6: exp_out = 32'h089351B3; // x = -2.7031, f(x) = 0.0670
          12'hEA7: exp_out = 32'h08A48989; // x = -2.6953, f(x) = 0.0675
          12'hEA8: exp_out = 32'h08B5E3F0; // x = -2.6875, f(x) = 0.0681
          12'hEA9: exp_out = 32'h08C76130; // x = -2.6797, f(x) = 0.0686
          12'hEAA: exp_out = 32'h08D9018C; // x = -2.6719, f(x) = 0.0691
          12'hEAB: exp_out = 32'h08EAC54D; // x = -2.6641, f(x) = 0.0697
          12'hEAC: exp_out = 32'h08FCACB9; // x = -2.6562, f(x) = 0.0702
          12'hEAD: exp_out = 32'h090EB818; // x = -2.6484, f(x) = 0.0708
          12'hEAE: exp_out = 32'h0920E7B2; // x = -2.6406, f(x) = 0.0713
          12'hEAF: exp_out = 32'h09333BCF; // x = -2.6328, f(x) = 0.0719
          12'hEB0: exp_out = 32'h0945B4BA; // x = -2.6250, f(x) = 0.0724
          12'hEB1: exp_out = 32'h095852BB; // x = -2.6172, f(x) = 0.0730
          12'hEB2: exp_out = 32'h096B161E; // x = -2.6094, f(x) = 0.0736
          12'hEB3: exp_out = 32'h097DFF2D; // x = -2.6016, f(x) = 0.0742
          12'hEB4: exp_out = 32'h09910E34; // x = -2.5938, f(x) = 0.0747
          12'hEB5: exp_out = 32'h09A4437F; // x = -2.5859, f(x) = 0.0753
          12'hEB6: exp_out = 32'h09B79F5B; // x = -2.5781, f(x) = 0.0759
          12'hEB7: exp_out = 32'h09CB2216; // x = -2.5703, f(x) = 0.0765
          12'hEB8: exp_out = 32'h09DECBFE; // x = -2.5625, f(x) = 0.0771
          12'hEB9: exp_out = 32'h09F29D60; // x = -2.5547, f(x) = 0.0777
          12'hEBA: exp_out = 32'h0A06968E; // x = -2.5469, f(x) = 0.0783
          12'hEBB: exp_out = 32'h0A1AB7D5; // x = -2.5391, f(x) = 0.0789
          12'hEBC: exp_out = 32'h0A2F0188; // x = -2.5312, f(x) = 0.0796
          12'hEBD: exp_out = 32'h0A4373F7; // x = -2.5234, f(x) = 0.0802
          12'hEBE: exp_out = 32'h0A580F73; // x = -2.5156, f(x) = 0.0808
          12'hEBF: exp_out = 32'h0A6CD450; // x = -2.5078, f(x) = 0.0814
          12'hEC0: exp_out = 32'h0A81C2E0; // x = -2.5000, f(x) = 0.0821
          12'hEC1: exp_out = 32'h0A96DB78; // x = -2.4922, f(x) = 0.0827
          12'hEC2: exp_out = 32'h0AAC1E6A; // x = -2.4844, f(x) = 0.0834
          12'hEC3: exp_out = 32'h0AC18C0E; // x = -2.4766, f(x) = 0.0840
          12'hEC4: exp_out = 32'h0AD724B7; // x = -2.4688, f(x) = 0.0847
          12'hEC5: exp_out = 32'h0AECE8BD; // x = -2.4609, f(x) = 0.0854
          12'hEC6: exp_out = 32'h0B02D877; // x = -2.4531, f(x) = 0.0860
          12'hEC7: exp_out = 32'h0B18F43D; // x = -2.4453, f(x) = 0.0867
          12'hEC8: exp_out = 32'h0B2F3C66; // x = -2.4375, f(x) = 0.0874
          12'hEC9: exp_out = 32'h0B45B14C; // x = -2.4297, f(x) = 0.0881
          12'hECA: exp_out = 32'h0B5C5349; // x = -2.4219, f(x) = 0.0888
          12'hECB: exp_out = 32'h0B7322B8; // x = -2.4141, f(x) = 0.0895
          12'hECC: exp_out = 32'h0B8A1FF3; // x = -2.4062, f(x) = 0.0902
          12'hECD: exp_out = 32'h0BA14B56; // x = -2.3984, f(x) = 0.0909
          12'hECE: exp_out = 32'h0BB8A53F; // x = -2.3906, f(x) = 0.0916
          12'hECF: exp_out = 32'h0BD02E0A; // x = -2.3828, f(x) = 0.0923
          12'hED0: exp_out = 32'h0BE7E617; // x = -2.3750, f(x) = 0.0930
          12'hED1: exp_out = 32'h0BFFCDC2; // x = -2.3672, f(x) = 0.0937
          12'hED2: exp_out = 32'h0C17E56E; // x = -2.3594, f(x) = 0.0945
          12'hED3: exp_out = 32'h0C302D78; // x = -2.3516, f(x) = 0.0952
          12'hED4: exp_out = 32'h0C48A644; // x = -2.3438, f(x) = 0.0960
          12'hED5: exp_out = 32'h0C615032; // x = -2.3359, f(x) = 0.0967
          12'hED6: exp_out = 32'h0C7A2BA6; // x = -2.3281, f(x) = 0.0975
          12'hED7: exp_out = 32'h0C933902; // x = -2.3203, f(x) = 0.0982
          12'hED8: exp_out = 32'h0CAC78AB; // x = -2.3125, f(x) = 0.0990
          12'hED9: exp_out = 32'h0CC5EB07; // x = -2.3047, f(x) = 0.0998
          12'hEDA: exp_out = 32'h0CDF907A; // x = -2.2969, f(x) = 0.1006
          12'hEDB: exp_out = 32'h0CF9696B; // x = -2.2891, f(x) = 0.1014
          12'hEDC: exp_out = 32'h0D137642; // x = -2.2812, f(x) = 0.1022
          12'hEDD: exp_out = 32'h0D2DB767; // x = -2.2734, f(x) = 0.1030
          12'hEDE: exp_out = 32'h0D482D43; // x = -2.2656, f(x) = 0.1038
          12'hEDF: exp_out = 32'h0D62D83F; // x = -2.2578, f(x) = 0.1046
          12'hEE0: exp_out = 32'h0D7DB8C7; // x = -2.2500, f(x) = 0.1054
          12'hEE1: exp_out = 32'h0D98CF46; // x = -2.2422, f(x) = 0.1062
          12'hEE2: exp_out = 32'h0DB41C29; // x = -2.2344, f(x) = 0.1071
          12'hEE3: exp_out = 32'h0DCF9FDB; // x = -2.2266, f(x) = 0.1079
          12'hEE4: exp_out = 32'h0DEB5ACD; // x = -2.2188, f(x) = 0.1087
          12'hEE5: exp_out = 32'h0E074D6C; // x = -2.2109, f(x) = 0.1096
          12'hEE6: exp_out = 32'h0E237828; // x = -2.2031, f(x) = 0.1105
          12'hEE7: exp_out = 32'h0E3FDB72; // x = -2.1953, f(x) = 0.1113
          12'hEE8: exp_out = 32'h0E5C77BC; // x = -2.1875, f(x) = 0.1122
          12'hEE9: exp_out = 32'h0E794D77; // x = -2.1797, f(x) = 0.1131
          12'hEEA: exp_out = 32'h0E965D18; // x = -2.1719, f(x) = 0.1140
          12'hEEB: exp_out = 32'h0EB3A713; // x = -2.1641, f(x) = 0.1149
          12'hEEC: exp_out = 32'h0ED12BDC; // x = -2.1562, f(x) = 0.1158
          12'hEED: exp_out = 32'h0EEEEBEA; // x = -2.1484, f(x) = 0.1167
          12'hEEE: exp_out = 32'h0F0CE7B3; // x = -2.1406, f(x) = 0.1176
          12'hEEF: exp_out = 32'h0F2B1FB0; // x = -2.1328, f(x) = 0.1185
          12'hEF0: exp_out = 32'h0F49945A; // x = -2.1250, f(x) = 0.1194
          12'hEF1: exp_out = 32'h0F68462B; // x = -2.1172, f(x) = 0.1204
          12'hEF2: exp_out = 32'h0F87359C; // x = -2.1094, f(x) = 0.1213
          12'hEF3: exp_out = 32'h0FA6632B; // x = -2.1016, f(x) = 0.1223
          12'hEF4: exp_out = 32'h0FC5CF53; // x = -2.0938, f(x) = 0.1232
          12'hEF5: exp_out = 32'h0FE57A92; // x = -2.0859, f(x) = 0.1242
          12'hEF6: exp_out = 32'h10056567; // x = -2.0781, f(x) = 0.1252
          12'hEF7: exp_out = 32'h10259052; // x = -2.0703, f(x) = 0.1261
          12'hEF8: exp_out = 32'h1045FBD4; // x = -2.0625, f(x) = 0.1271
          12'hEF9: exp_out = 32'h1066A86D; // x = -2.0547, f(x) = 0.1281
          12'hEFA: exp_out = 32'h108796A1; // x = -2.0469, f(x) = 0.1291
          12'hEFB: exp_out = 32'h10A8C6F4; // x = -2.0391, f(x) = 0.1302
          12'hEFC: exp_out = 32'h10CA39E9; // x = -2.0312, f(x) = 0.1312
          12'hEFD: exp_out = 32'h10EBF008; // x = -2.0234, f(x) = 0.1322
          12'hEFE: exp_out = 32'h110DE9D6; // x = -2.0156, f(x) = 0.1332
          12'hEFF: exp_out = 32'h113027DD; // x = -2.0078, f(x) = 0.1343
          12'hF00: exp_out = 32'h1152AAA4; // x = -2.0000, f(x) = 0.1353
          12'hF01: exp_out = 32'h117572B6; // x = -1.9922, f(x) = 0.1364
          12'hF02: exp_out = 32'h1198809D; // x = -1.9844, f(x) = 0.1375
          12'hF03: exp_out = 32'h11BBD4E7; // x = -1.9766, f(x) = 0.1385
          12'hF04: exp_out = 32'h11DF7020; // x = -1.9688, f(x) = 0.1396
          12'hF05: exp_out = 32'h120352D7; // x = -1.9609, f(x) = 0.1407
          12'hF06: exp_out = 32'h12277D9B; // x = -1.9531, f(x) = 0.1418
          12'hF07: exp_out = 32'h124BF0FE; // x = -1.9453, f(x) = 0.1429
          12'hF08: exp_out = 32'h1270AD90; // x = -1.9375, f(x) = 0.1441
          12'hF09: exp_out = 32'h1295B3E5; // x = -1.9297, f(x) = 0.1452
          12'hF0A: exp_out = 32'h12BB0491; // x = -1.9219, f(x) = 0.1463
          12'hF0B: exp_out = 32'h12E0A02A; // x = -1.9141, f(x) = 0.1475
          12'hF0C: exp_out = 32'h13068744; // x = -1.9062, f(x) = 0.1486
          12'hF0D: exp_out = 32'h132CBA79; // x = -1.8984, f(x) = 0.1498
          12'hF0E: exp_out = 32'h13533A61; // x = -1.8906, f(x) = 0.1510
          12'hF0F: exp_out = 32'h137A0796; // x = -1.8828, f(x) = 0.1522
          12'hF10: exp_out = 32'h13A122B4; // x = -1.8750, f(x) = 0.1534
          12'hF11: exp_out = 32'h13C88C56; // x = -1.8672, f(x) = 0.1546
          12'hF12: exp_out = 32'h13F0451A; // x = -1.8594, f(x) = 0.1558
          12'hF13: exp_out = 32'h14184D9F; // x = -1.8516, f(x) = 0.1570
          12'hF14: exp_out = 32'h1440A686; // x = -1.8438, f(x) = 0.1582
          12'hF15: exp_out = 32'h1469506F; // x = -1.8359, f(x) = 0.1595
          12'hF16: exp_out = 32'h14924BFE; // x = -1.8281, f(x) = 0.1607
          12'hF17: exp_out = 32'h14BB99D6; // x = -1.8203, f(x) = 0.1620
          12'hF18: exp_out = 32'h14E53A9D; // x = -1.8125, f(x) = 0.1632
          12'hF19: exp_out = 32'h150F2EF8; // x = -1.8047, f(x) = 0.1645
          12'hF1A: exp_out = 32'h15397791; // x = -1.7969, f(x) = 0.1658
          12'hF1B: exp_out = 32'h1564150F; // x = -1.7891, f(x) = 0.1671
          12'hF1C: exp_out = 32'h158F081E; // x = -1.7812, f(x) = 0.1684
          12'hF1D: exp_out = 32'h15BA5169; // x = -1.7734, f(x) = 0.1697
          12'hF1E: exp_out = 32'h15E5F19E; // x = -1.7656, f(x) = 0.1711
          12'hF1F: exp_out = 32'h1611E96A; // x = -1.7578, f(x) = 0.1724
          12'hF20: exp_out = 32'h163E397E; // x = -1.7500, f(x) = 0.1738
          12'hF21: exp_out = 32'h166AE28B; // x = -1.7422, f(x) = 0.1751
          12'hF22: exp_out = 32'h1697E544; // x = -1.7344, f(x) = 0.1765
          12'hF23: exp_out = 32'h16C5425C; // x = -1.7266, f(x) = 0.1779
          12'hF24: exp_out = 32'h16F2FA8A; // x = -1.7188, f(x) = 0.1793
          12'hF25: exp_out = 32'h17210E84; // x = -1.7109, f(x) = 0.1807
          12'hF26: exp_out = 32'h174F7F02; // x = -1.7031, f(x) = 0.1821
          12'hF27: exp_out = 32'h177E4CBE; // x = -1.6953, f(x) = 0.1835
          12'hF28: exp_out = 32'h17AD7873; // x = -1.6875, f(x) = 0.1850
          12'hF29: exp_out = 32'h17DD02DF; // x = -1.6797, f(x) = 0.1864
          12'hF2A: exp_out = 32'h180CECBF; // x = -1.6719, f(x) = 0.1879
          12'hF2B: exp_out = 32'h183D36D2; // x = -1.6641, f(x) = 0.1894
          12'hF2C: exp_out = 32'h186DE1DB; // x = -1.6562, f(x) = 0.1909
          12'hF2D: exp_out = 32'h189EEE9B; // x = -1.6484, f(x) = 0.1924
          12'hF2E: exp_out = 32'h18D05DD7; // x = -1.6406, f(x) = 0.1939
          12'hF2F: exp_out = 32'h19023054; // x = -1.6328, f(x) = 0.1954
          12'hF30: exp_out = 32'h193466DB; // x = -1.6250, f(x) = 0.1969
          12'hF31: exp_out = 32'h19670233; // x = -1.6172, f(x) = 0.1985
          12'hF32: exp_out = 32'h199A0327; // x = -1.6094, f(x) = 0.2000
          12'hF33: exp_out = 32'h19CD6A84; // x = -1.6016, f(x) = 0.2016
          12'hF34: exp_out = 32'h1A013916; // x = -1.5938, f(x) = 0.2032
          12'hF35: exp_out = 32'h1A356FAD; // x = -1.5859, f(x) = 0.2048
          12'hF36: exp_out = 32'h1A6A0F1B; // x = -1.5781, f(x) = 0.2064
          12'hF37: exp_out = 32'h1A9F1830; // x = -1.5703, f(x) = 0.2080
          12'hF38: exp_out = 32'h1AD48BC2; // x = -1.5625, f(x) = 0.2096
          12'hF39: exp_out = 32'h1B0A6AA7; // x = -1.5547, f(x) = 0.2113
          12'hF3A: exp_out = 32'h1B40B5B5; // x = -1.5469, f(x) = 0.2129
          12'hF3B: exp_out = 32'h1B776DC6; // x = -1.5391, f(x) = 0.2146
          12'hF3C: exp_out = 32'h1BAE93B5; // x = -1.5312, f(x) = 0.2163
          12'hF3D: exp_out = 32'h1BE6285F; // x = -1.5234, f(x) = 0.2180
          12'hF3E: exp_out = 32'h1C1E2CA1; // x = -1.5156, f(x) = 0.2197
          12'hF3F: exp_out = 32'h1C56A15C; // x = -1.5078, f(x) = 0.2214
          12'hF40: exp_out = 32'h1C8F8772; // x = -1.5000, f(x) = 0.2231
          12'hF41: exp_out = 32'h1CC8DFC6; // x = -1.4922, f(x) = 0.2249
          12'hF42: exp_out = 32'h1D02AB3E; // x = -1.4844, f(x) = 0.2266
          12'hF43: exp_out = 32'h1D3CEAC1; // x = -1.4766, f(x) = 0.2284
          12'hF44: exp_out = 32'h1D779F37; // x = -1.4688, f(x) = 0.2302
          12'hF45: exp_out = 32'h1DB2C98C; // x = -1.4609, f(x) = 0.2320
          12'hF46: exp_out = 32'h1DEE6AAD; // x = -1.4531, f(x) = 0.2338
          12'hF47: exp_out = 32'h1E2A8387; // x = -1.4453, f(x) = 0.2357
          12'hF48: exp_out = 32'h1E67150B; // x = -1.4375, f(x) = 0.2375
          12'hF49: exp_out = 32'h1EA4202C; // x = -1.4297, f(x) = 0.2394
          12'hF4A: exp_out = 32'h1EE1A5DD; // x = -1.4219, f(x) = 0.2413
          12'hF4B: exp_out = 32'h1F1FA716; // x = -1.4141, f(x) = 0.2432
          12'hF4C: exp_out = 32'h1F5E24CD; // x = -1.4062, f(x) = 0.2451
          12'hF4D: exp_out = 32'h1F9D1FFD; // x = -1.3984, f(x) = 0.2470
          12'hF4E: exp_out = 32'h1FDC99A1; // x = -1.3906, f(x) = 0.2489
          12'hF4F: exp_out = 32'h201C92B8; // x = -1.3828, f(x) = 0.2509
          12'hF50: exp_out = 32'h205D0C42; // x = -1.3750, f(x) = 0.2528
          12'hF51: exp_out = 32'h209E073F; // x = -1.3672, f(x) = 0.2548
          12'hF52: exp_out = 32'h20DF84B6; // x = -1.3594, f(x) = 0.2568
          12'hF53: exp_out = 32'h212185AA; // x = -1.3516, f(x) = 0.2588
          12'hF54: exp_out = 32'h21640B25; // x = -1.3438, f(x) = 0.2609
          12'hF55: exp_out = 32'h21A71630; // x = -1.3359, f(x) = 0.2629
          12'hF56: exp_out = 32'h21EAA7D7; // x = -1.3281, f(x) = 0.2650
          12'hF57: exp_out = 32'h222EC129; // x = -1.3203, f(x) = 0.2671
          12'hF58: exp_out = 32'h22736337; // x = -1.3125, f(x) = 0.2691
          12'hF59: exp_out = 32'h22B88F12; // x = -1.3047, f(x) = 0.2713
          12'hF5A: exp_out = 32'h22FE45D0; // x = -1.2969, f(x) = 0.2734
          12'hF5B: exp_out = 32'h23448887; // x = -1.2891, f(x) = 0.2755
          12'hF5C: exp_out = 32'h238B5850; // x = -1.2812, f(x) = 0.2777
          12'hF5D: exp_out = 32'h23D2B647; // x = -1.2734, f(x) = 0.2799
          12'hF5E: exp_out = 32'h241AA388; // x = -1.2656, f(x) = 0.2821
          12'hF5F: exp_out = 32'h24632135; // x = -1.2578, f(x) = 0.2843
          12'hF60: exp_out = 32'h24AC306E; // x = -1.2500, f(x) = 0.2865
          12'hF61: exp_out = 32'h24F5D259; // x = -1.2422, f(x) = 0.2888
          12'hF62: exp_out = 32'h2540081A; // x = -1.2344, f(x) = 0.2910
          12'hF63: exp_out = 32'h258AD2DC; // x = -1.2266, f(x) = 0.2933
          12'hF64: exp_out = 32'h25D633CA; // x = -1.2188, f(x) = 0.2956
          12'hF65: exp_out = 32'h26222C10; // x = -1.2109, f(x) = 0.2979
          12'hF66: exp_out = 32'h266EBCE0; // x = -1.2031, f(x) = 0.3003
          12'hF67: exp_out = 32'h26BBE76A; // x = -1.1953, f(x) = 0.3026
          12'hF68: exp_out = 32'h2709ACE5; // x = -1.1875, f(x) = 0.3050
          12'hF69: exp_out = 32'h27580E86; // x = -1.1797, f(x) = 0.3074
          12'hF6A: exp_out = 32'h27A70D88; // x = -1.1719, f(x) = 0.3098
          12'hF6B: exp_out = 32'h27F6AB26; // x = -1.1641, f(x) = 0.3122
          12'hF6C: exp_out = 32'h2846E89F; // x = -1.1562, f(x) = 0.3147
          12'hF6D: exp_out = 32'h2897C734; // x = -1.1484, f(x) = 0.3171
          12'hF6E: exp_out = 32'h28E94828; // x = -1.1406, f(x) = 0.3196
          12'hF6F: exp_out = 32'h293B6CC1; // x = -1.1328, f(x) = 0.3221
          12'hF70: exp_out = 32'h298E3649; // x = -1.1250, f(x) = 0.3247
          12'hF71: exp_out = 32'h29E1A609; // x = -1.1172, f(x) = 0.3272
          12'hF72: exp_out = 32'h2A35BD51; // x = -1.1094, f(x) = 0.3298
          12'hF73: exp_out = 32'h2A8A7D6F; // x = -1.1016, f(x) = 0.3324
          12'hF74: exp_out = 32'h2ADFE7B8; // x = -1.0938, f(x) = 0.3350
          12'hF75: exp_out = 32'h2B35FD80; // x = -1.0859, f(x) = 0.3376
          12'hF76: exp_out = 32'h2B8CC021; // x = -1.0781, f(x) = 0.3402
          12'hF77: exp_out = 32'h2BE430F5; // x = -1.0703, f(x) = 0.3429
          12'hF78: exp_out = 32'h2C3C515A; // x = -1.0625, f(x) = 0.3456
          12'hF79: exp_out = 32'h2C9522B0; // x = -1.0547, f(x) = 0.3483
          12'hF7A: exp_out = 32'h2CEEA65C; // x = -1.0469, f(x) = 0.3510
          12'hF7B: exp_out = 32'h2D48DDC2; // x = -1.0391, f(x) = 0.3538
          12'hF7C: exp_out = 32'h2DA3CA4B; // x = -1.0312, f(x) = 0.3566
          12'hF7D: exp_out = 32'h2DFF6D65; // x = -1.0234, f(x) = 0.3594
          12'hF7E: exp_out = 32'h2E5BC87C; // x = -1.0156, f(x) = 0.3622
          12'hF7F: exp_out = 32'h2EB8DD02; // x = -1.0078, f(x) = 0.3650
          12'hF80: exp_out = 32'h2F16AC6C; // x = -1.0000, f(x) = 0.3679
          12'hF81: exp_out = 32'h2F753831; // x = -0.9922, f(x) = 0.3708
          12'hF82: exp_out = 32'h2FD481CC; // x = -0.9844, f(x) = 0.3737
          12'hF83: exp_out = 32'h30348AB8; // x = -0.9766, f(x) = 0.3766
          12'hF84: exp_out = 32'h30955477; // x = -0.9688, f(x) = 0.3796
          12'hF85: exp_out = 32'h30F6E08C; // x = -0.9609, f(x) = 0.3825
          12'hF86: exp_out = 32'h3159307C; // x = -0.9531, f(x) = 0.3855
          12'hF87: exp_out = 32'h31BC45D1; // x = -0.9453, f(x) = 0.3886
          12'hF88: exp_out = 32'h32202218; // x = -0.9375, f(x) = 0.3916
          12'hF89: exp_out = 32'h3284C6DF; // x = -0.9297, f(x) = 0.3947
          12'hF8A: exp_out = 32'h32EA35BA; // x = -0.9219, f(x) = 0.3978
          12'hF8B: exp_out = 32'h3350703E; // x = -0.9141, f(x) = 0.4009
          12'hF8C: exp_out = 32'h33B77804; // x = -0.9062, f(x) = 0.4040
          12'hF8D: exp_out = 32'h341F4EA8; // x = -0.8984, f(x) = 0.4072
          12'hF8E: exp_out = 32'h3487F5C9; // x = -0.8906, f(x) = 0.4104
          12'hF8F: exp_out = 32'h34F16F0B; // x = -0.8828, f(x) = 0.4136
          12'hF90: exp_out = 32'h355BBC13; // x = -0.8750, f(x) = 0.4169
          12'hF91: exp_out = 32'h35C6DE8A; // x = -0.8672, f(x) = 0.4201
          12'hF92: exp_out = 32'h3632D81C; // x = -0.8594, f(x) = 0.4234
          12'hF93: exp_out = 32'h369FAA7B; // x = -0.8516, f(x) = 0.4267
          12'hF94: exp_out = 32'h370D5758; // x = -0.8438, f(x) = 0.4301
          12'hF95: exp_out = 32'h377BE06B; // x = -0.8359, f(x) = 0.4335
          12'hF96: exp_out = 32'h37EB476D; // x = -0.8281, f(x) = 0.4369
          12'hF97: exp_out = 32'h385B8E1E; // x = -0.8203, f(x) = 0.4403
          12'hF98: exp_out = 32'h38CCB63C; // x = -0.8125, f(x) = 0.4437
          12'hF99: exp_out = 32'h393EC18E; // x = -0.8047, f(x) = 0.4472
          12'hF9A: exp_out = 32'h39B1B1DB; // x = -0.7969, f(x) = 0.4507
          12'hF9B: exp_out = 32'h3A2588EF; // x = -0.7891, f(x) = 0.4543
          12'hF9C: exp_out = 32'h3A9A489A; // x = -0.7812, f(x) = 0.4578
          12'hF9D: exp_out = 32'h3B0FF2AE; // x = -0.7734, f(x) = 0.4614
          12'hF9E: exp_out = 32'h3B868902; // x = -0.7656, f(x) = 0.4650
          12'hF9F: exp_out = 32'h3BFE0D71; // x = -0.7578, f(x) = 0.4687
          12'hFA0: exp_out = 32'h3C7681D8; // x = -0.7500, f(x) = 0.4724
          12'hFA1: exp_out = 32'h3CEFE819; // x = -0.7422, f(x) = 0.4761
          12'hFA2: exp_out = 32'h3D6A421B; // x = -0.7344, f(x) = 0.4798
          12'hFA3: exp_out = 32'h3DE591C6; // x = -0.7266, f(x) = 0.4836
          12'hFA4: exp_out = 32'h3E61D907; // x = -0.7188, f(x) = 0.4874
          12'hFA5: exp_out = 32'h3EDF19D0; // x = -0.7109, f(x) = 0.4912
          12'hFA6: exp_out = 32'h3F5D5616; // x = -0.7031, f(x) = 0.4950
          12'hFA7: exp_out = 32'h3FDC8FD1; // x = -0.6953, f(x) = 0.4989
          12'hFA8: exp_out = 32'h405CC8FF; // x = -0.6875, f(x) = 0.5028
          12'hFA9: exp_out = 32'h40DE03A1; // x = -0.6797, f(x) = 0.5068
          12'hFAA: exp_out = 32'h416041BB; // x = -0.6719, f(x) = 0.5108
          12'hFAB: exp_out = 32'h41E38556; // x = -0.6641, f(x) = 0.5148
          12'hFAC: exp_out = 32'h4267D080; // x = -0.6562, f(x) = 0.5188
          12'hFAD: exp_out = 32'h42ED2549; // x = -0.6484, f(x) = 0.5229
          12'hFAE: exp_out = 32'h437385C8; // x = -0.6406, f(x) = 0.5270
          12'hFAF: exp_out = 32'h43FAF414; // x = -0.6328, f(x) = 0.5311
          12'hFB0: exp_out = 32'h4483724D; // x = -0.6250, f(x) = 0.5353
          12'hFB1: exp_out = 32'h450D0294; // x = -0.6172, f(x) = 0.5395
          12'hFB2: exp_out = 32'h4597A710; // x = -0.6094, f(x) = 0.5437
          12'hFB3: exp_out = 32'h462361EA; // x = -0.6016, f(x) = 0.5480
          12'hFB4: exp_out = 32'h46B03552; // x = -0.5938, f(x) = 0.5523
          12'hFB5: exp_out = 32'h473E237C; // x = -0.5859, f(x) = 0.5566
          12'hFB6: exp_out = 32'h47CD2E9E; // x = -0.5781, f(x) = 0.5609
          12'hFB7: exp_out = 32'h485D58F6; // x = -0.5703, f(x) = 0.5653
          12'hFB8: exp_out = 32'h48EEA4C3; // x = -0.5625, f(x) = 0.5698
          12'hFB9: exp_out = 32'h4981144B; // x = -0.5547, f(x) = 0.5743
          12'hFBA: exp_out = 32'h4A14A9D8; // x = -0.5469, f(x) = 0.5788
          12'hFBB: exp_out = 32'h4AA967B8; // x = -0.5391, f(x) = 0.5833
          12'hFBC: exp_out = 32'h4B3F503E; // x = -0.5312, f(x) = 0.5879
          12'hFBD: exp_out = 32'h4BD665C2; // x = -0.5234, f(x) = 0.5925
          12'hFBE: exp_out = 32'h4C6EAA9F; // x = -0.5156, f(x) = 0.5971
          12'hFBF: exp_out = 32'h4D082138; // x = -0.5078, f(x) = 0.6018
          12'hFC0: exp_out = 32'h4DA2CBF2; // x = -0.5000, f(x) = 0.6065
          12'hFC1: exp_out = 32'h4E3EAD37; // x = -0.4922, f(x) = 0.6113
          12'hFC2: exp_out = 32'h4EDBC777; // x = -0.4844, f(x) = 0.6161
          12'hFC3: exp_out = 32'h4F7A1D27; // x = -0.4766, f(x) = 0.6209
          12'hFC4: exp_out = 32'h5019B0C0; // x = -0.4688, f(x) = 0.6258
          12'hFC5: exp_out = 32'h50BA84C0; // x = -0.4609, f(x) = 0.6307
          12'hFC6: exp_out = 32'h515C9BAA; // x = -0.4531, f(x) = 0.6356
          12'hFC7: exp_out = 32'h51FFF807; // x = -0.4453, f(x) = 0.6406
          12'hFC8: exp_out = 32'h52A49C65; // x = -0.4375, f(x) = 0.6456
          12'hFC9: exp_out = 32'h534A8B55; // x = -0.4297, f(x) = 0.6507
          12'hFCA: exp_out = 32'h53F1C770; // x = -0.4219, f(x) = 0.6558
          12'hFCB: exp_out = 32'h549A5353; // x = -0.4141, f(x) = 0.6610
          12'hFCC: exp_out = 32'h5544319F; // x = -0.4062, f(x) = 0.6661
          12'hFCD: exp_out = 32'h55EF64FD; // x = -0.3984, f(x) = 0.6714
          12'hFCE: exp_out = 32'h569BF018; // x = -0.3906, f(x) = 0.6766
          12'hFCF: exp_out = 32'h5749D5A4; // x = -0.3828, f(x) = 0.6819
          12'hFD0: exp_out = 32'h57F91858; // x = -0.3750, f(x) = 0.6873
          12'hFD1: exp_out = 32'h58A9BAF0; // x = -0.3672, f(x) = 0.6927
          12'hFD2: exp_out = 32'h595BC030; // x = -0.3594, f(x) = 0.6981
          12'hFD3: exp_out = 32'h5A0F2ADF; // x = -0.3516, f(x) = 0.7036
          12'hFD4: exp_out = 32'h5AC3FDCB; // x = -0.3438, f(x) = 0.7091
          12'hFD5: exp_out = 32'h5B7A3BC8; // x = -0.3359, f(x) = 0.7147
          12'hFD6: exp_out = 32'h5C31E7AF; // x = -0.3281, f(x) = 0.7203
          12'hFD7: exp_out = 32'h5CEB045D; // x = -0.3203, f(x) = 0.7259
          12'hFD8: exp_out = 32'h5DA594B8; // x = -0.3125, f(x) = 0.7316
          12'hFD9: exp_out = 32'h5E619BA9; // x = -0.3047, f(x) = 0.7374
          12'hFDA: exp_out = 32'h5F1F1C22; // x = -0.2969, f(x) = 0.7431
          12'hFDB: exp_out = 32'h5FDE1918; // x = -0.2891, f(x) = 0.7490
          12'hFDC: exp_out = 32'h609E9586; // x = -0.2812, f(x) = 0.7548
          12'hFDD: exp_out = 32'h6160946F; // x = -0.2734, f(x) = 0.7608
          12'hFDE: exp_out = 32'h622418DC; // x = -0.2656, f(x) = 0.7667
          12'hFDF: exp_out = 32'h62E925D9; // x = -0.2578, f(x) = 0.7727
          12'hFE0: exp_out = 32'h63AFBE7B; // x = -0.2500, f(x) = 0.7788
          12'hFE1: exp_out = 32'h6477E5DC; // x = -0.2422, f(x) = 0.7849
          12'hFE2: exp_out = 32'h65419F1E; // x = -0.2344, f(x) = 0.7911
          12'hFE3: exp_out = 32'h660CED67; // x = -0.2266, f(x) = 0.7973
          12'hFE4: exp_out = 32'h66D9D3E4; // x = -0.2188, f(x) = 0.8035
          12'hFE5: exp_out = 32'h67A855C9; // x = -0.2109, f(x) = 0.8098
          12'hFE6: exp_out = 32'h6878764F; // x = -0.2031, f(x) = 0.8162
          12'hFE7: exp_out = 32'h694A38B8; // x = -0.1953, f(x) = 0.8226
          12'hFE8: exp_out = 32'h6A1DA04B; // x = -0.1875, f(x) = 0.8290
          12'hFE9: exp_out = 32'h6AF2B055; // x = -0.1797, f(x) = 0.8355
          12'hFEA: exp_out = 32'h6BC96C2A; // x = -0.1719, f(x) = 0.8421
          12'hFEB: exp_out = 32'h6CA1D725; // x = -0.1641, f(x) = 0.8487
          12'hFEC: exp_out = 32'h6D7BF4A8; // x = -0.1562, f(x) = 0.8553
          12'hFED: exp_out = 32'h6E57C81B; // x = -0.1484, f(x) = 0.8621
          12'hFEE: exp_out = 32'h6F3554EE; // x = -0.1406, f(x) = 0.8688
          12'hFEF: exp_out = 32'h70149E98; // x = -0.1328, f(x) = 0.8756
          12'hFF0: exp_out = 32'h70F5A894; // x = -0.1250, f(x) = 0.8825
          12'hFF1: exp_out = 32'h71D87667; // x = -0.1172, f(x) = 0.8894
          12'hFF2: exp_out = 32'h72BD0B9D; // x = -0.1094, f(x) = 0.8964
          12'hFF3: exp_out = 32'h73A36BC8; // x = -0.1016, f(x) = 0.9034
          12'hFF4: exp_out = 32'h748B9A80; // x = -0.0938, f(x) = 0.9105
          12'hFF5: exp_out = 32'h75759B68; // x = -0.0859, f(x) = 0.9177
          12'hFF6: exp_out = 32'h76617227; // x = -0.0781, f(x) = 0.9248
          12'hFF7: exp_out = 32'h774F226D; // x = -0.0703, f(x) = 0.9321
          12'hFF8: exp_out = 32'h783EAFEF; // x = -0.0625, f(x) = 0.9394
          12'hFF9: exp_out = 32'h79301E6D; // x = -0.0547, f(x) = 0.9468
          12'hFFA: exp_out = 32'h7A2371AC; // x = -0.0469, f(x) = 0.9542
          12'hFFB: exp_out = 32'h7B18AD79; // x = -0.0391, f(x) = 0.9617
          12'hFFC: exp_out = 32'h7C0FD5AA; // x = -0.0312, f(x) = 0.9692
          12'hFFD: exp_out = 32'h7D08EE1B; // x = -0.0234, f(x) = 0.9768
          12'hFFE: exp_out = 32'h7E03FAB0; // x = -0.0156, f(x) = 0.9845
          12'hFFF: exp_out = 32'h7F00FF56; // x = -0.0078, f(x) = 0.9922
          default: exp_out = 32'h0; 
        endcase
end

wire [11:0] soft_addr = input_data0[31:20];
reg  [31:0] soft_out;
always @( * ) begin
  case ( soft_addr )
    12'h000: soft_out = 32'h7FFFFFFF; 
    12'h800: soft_out = 32'h00000000; // x = -32.0000, f(x) = 0.0000
    12'h801: soft_out = 32'h00000000; // x = -31.9844, f(x) = 0.0000
    12'h802: soft_out = 32'h00000000; // x = -31.9688, f(x) = 0.0000
    12'h803: soft_out = 32'h00000000; // x = -31.9531, f(x) = 0.0000
    12'h804: soft_out = 32'h00000000; // x = -31.9375, f(x) = 0.0000
    12'h805: soft_out = 32'h00000000; // x = -31.9219, f(x) = 0.0000
    12'h806: soft_out = 32'h00000000; // x = -31.9062, f(x) = 0.0000
    12'h807: soft_out = 32'h00000000; // x = -31.8906, f(x) = 0.0000
    12'h808: soft_out = 32'h00000000; // x = -31.8750, f(x) = 0.0000
    12'h809: soft_out = 32'h00000000; // x = -31.8594, f(x) = 0.0000
    12'h80A: soft_out = 32'h00000000; // x = -31.8438, f(x) = 0.0000
    12'h80B: soft_out = 32'h00000000; // x = -31.8281, f(x) = 0.0000
    12'h80C: soft_out = 32'h00000000; // x = -31.8125, f(x) = 0.0000
    12'h80D: soft_out = 32'h00000000; // x = -31.7969, f(x) = 0.0000
    12'h80E: soft_out = 32'h00000000; // x = -31.7812, f(x) = 0.0000
    12'h80F: soft_out = 32'h00000000; // x = -31.7656, f(x) = 0.0000
    12'h810: soft_out = 32'h00000000; // x = -31.7500, f(x) = 0.0000
    12'h811: soft_out = 32'h00000000; // x = -31.7344, f(x) = 0.0000
    12'h812: soft_out = 32'h00000000; // x = -31.7188, f(x) = 0.0000
    12'h813: soft_out = 32'h00000000; // x = -31.7031, f(x) = 0.0000
    12'h814: soft_out = 32'h00000000; // x = -31.6875, f(x) = 0.0000
    12'h815: soft_out = 32'h00000000; // x = -31.6719, f(x) = 0.0000
    12'h816: soft_out = 32'h00000000; // x = -31.6562, f(x) = 0.0000
    12'h817: soft_out = 32'h00000000; // x = -31.6406, f(x) = 0.0000
    12'h818: soft_out = 32'h00000000; // x = -31.6250, f(x) = 0.0000
    12'h819: soft_out = 32'h00000000; // x = -31.6094, f(x) = 0.0000
    12'h81A: soft_out = 32'h00000000; // x = -31.5938, f(x) = 0.0000
    12'h81B: soft_out = 32'h00000000; // x = -31.5781, f(x) = 0.0000
    12'h81C: soft_out = 32'h00000000; // x = -31.5625, f(x) = 0.0000
    12'h81D: soft_out = 32'h00000000; // x = -31.5469, f(x) = 0.0000
    12'h81E: soft_out = 32'h00000000; // x = -31.5312, f(x) = 0.0000
    12'h81F: soft_out = 32'h00000000; // x = -31.5156, f(x) = 0.0000
    12'h820: soft_out = 32'h00000000; // x = -31.5000, f(x) = 0.0000
    12'h821: soft_out = 32'h00000000; // x = -31.4844, f(x) = 0.0000
    12'h822: soft_out = 32'h00000000; // x = -31.4688, f(x) = 0.0000
    12'h823: soft_out = 32'h00000000; // x = -31.4531, f(x) = 0.0000
    12'h824: soft_out = 32'h00000000; // x = -31.4375, f(x) = 0.0000
    12'h825: soft_out = 32'h00000000; // x = -31.4219, f(x) = 0.0000
    12'h826: soft_out = 32'h00000000; // x = -31.4062, f(x) = 0.0000
    12'h827: soft_out = 32'h00000000; // x = -31.3906, f(x) = 0.0000
    12'h828: soft_out = 32'h00000000; // x = -31.3750, f(x) = 0.0000
    12'h829: soft_out = 32'h00000000; // x = -31.3594, f(x) = 0.0000
    12'h82A: soft_out = 32'h00000000; // x = -31.3438, f(x) = 0.0000
    12'h82B: soft_out = 32'h00000000; // x = -31.3281, f(x) = 0.0000
    12'h82C: soft_out = 32'h00000000; // x = -31.3125, f(x) = 0.0000
    12'h82D: soft_out = 32'h00000000; // x = -31.2969, f(x) = 0.0000
    12'h82E: soft_out = 32'h00000000; // x = -31.2812, f(x) = 0.0000
    12'h82F: soft_out = 32'h00000000; // x = -31.2656, f(x) = 0.0000
    12'h830: soft_out = 32'h00000000; // x = -31.2500, f(x) = 0.0000
    12'h831: soft_out = 32'h00000000; // x = -31.2344, f(x) = 0.0000
    12'h832: soft_out = 32'h00000000; // x = -31.2188, f(x) = 0.0000
    12'h833: soft_out = 32'h00000000; // x = -31.2031, f(x) = 0.0000
    12'h834: soft_out = 32'h00000000; // x = -31.1875, f(x) = 0.0000
    12'h835: soft_out = 32'h00000000; // x = -31.1719, f(x) = 0.0000
    12'h836: soft_out = 32'h00000000; // x = -31.1562, f(x) = 0.0000
    12'h837: soft_out = 32'h00000000; // x = -31.1406, f(x) = 0.0000
    12'h838: soft_out = 32'h00000000; // x = -31.1250, f(x) = 0.0000
    12'h839: soft_out = 32'h00000000; // x = -31.1094, f(x) = 0.0000
    12'h83A: soft_out = 32'h00000000; // x = -31.0938, f(x) = 0.0000
    12'h83B: soft_out = 32'h00000000; // x = -31.0781, f(x) = 0.0000
    12'h83C: soft_out = 32'h00000000; // x = -31.0625, f(x) = 0.0000
    12'h83D: soft_out = 32'h00000000; // x = -31.0469, f(x) = 0.0000
    12'h83E: soft_out = 32'h00000000; // x = -31.0312, f(x) = 0.0000
    12'h83F: soft_out = 32'h00000000; // x = -31.0156, f(x) = 0.0000
    12'h840: soft_out = 32'h00000000; // x = -31.0000, f(x) = 0.0000
    12'h841: soft_out = 32'h00000000; // x = -30.9844, f(x) = 0.0000
    12'h842: soft_out = 32'h00000000; // x = -30.9688, f(x) = 0.0000
    12'h843: soft_out = 32'h00000000; // x = -30.9531, f(x) = 0.0000
    12'h844: soft_out = 32'h00000000; // x = -30.9375, f(x) = 0.0000
    12'h845: soft_out = 32'h00000000; // x = -30.9219, f(x) = 0.0000
    12'h846: soft_out = 32'h00000000; // x = -30.9062, f(x) = 0.0000
    12'h847: soft_out = 32'h00000000; // x = -30.8906, f(x) = 0.0000
    12'h848: soft_out = 32'h00000000; // x = -30.8750, f(x) = 0.0000
    12'h849: soft_out = 32'h00000000; // x = -30.8594, f(x) = 0.0000
    12'h84A: soft_out = 32'h00000000; // x = -30.8438, f(x) = 0.0000
    12'h84B: soft_out = 32'h00000000; // x = -30.8281, f(x) = 0.0000
    12'h84C: soft_out = 32'h00000000; // x = -30.8125, f(x) = 0.0000
    12'h84D: soft_out = 32'h00000000; // x = -30.7969, f(x) = 0.0000
    12'h84E: soft_out = 32'h00000000; // x = -30.7812, f(x) = 0.0000
    12'h84F: soft_out = 32'h00000000; // x = -30.7656, f(x) = 0.0000
    12'h850: soft_out = 32'h00000000; // x = -30.7500, f(x) = 0.0000
    12'h851: soft_out = 32'h00000000; // x = -30.7344, f(x) = 0.0000
    12'h852: soft_out = 32'h00000000; // x = -30.7188, f(x) = 0.0000
    12'h853: soft_out = 32'h00000000; // x = -30.7031, f(x) = 0.0000
    12'h854: soft_out = 32'h00000000; // x = -30.6875, f(x) = 0.0000
    12'h855: soft_out = 32'h00000000; // x = -30.6719, f(x) = 0.0000
    12'h856: soft_out = 32'h00000000; // x = -30.6562, f(x) = 0.0000
    12'h857: soft_out = 32'h00000000; // x = -30.6406, f(x) = 0.0000
    12'h858: soft_out = 32'h00000000; // x = -30.6250, f(x) = 0.0000
    12'h859: soft_out = 32'h00000000; // x = -30.6094, f(x) = 0.0000
    12'h85A: soft_out = 32'h00000000; // x = -30.5938, f(x) = 0.0000
    12'h85B: soft_out = 32'h00000000; // x = -30.5781, f(x) = 0.0000
    12'h85C: soft_out = 32'h00000000; // x = -30.5625, f(x) = 0.0000
    12'h85D: soft_out = 32'h00000000; // x = -30.5469, f(x) = 0.0000
    12'h85E: soft_out = 32'h00000000; // x = -30.5312, f(x) = 0.0000
    12'h85F: soft_out = 32'h00000000; // x = -30.5156, f(x) = 0.0000
    12'h860: soft_out = 32'h00000000; // x = -30.5000, f(x) = 0.0000
    12'h861: soft_out = 32'h00000000; // x = -30.4844, f(x) = 0.0000
    12'h862: soft_out = 32'h00000000; // x = -30.4688, f(x) = 0.0000
    12'h863: soft_out = 32'h00000000; // x = -30.4531, f(x) = 0.0000
    12'h864: soft_out = 32'h00000000; // x = -30.4375, f(x) = 0.0000
    12'h865: soft_out = 32'h00000000; // x = -30.4219, f(x) = 0.0000
    12'h866: soft_out = 32'h00000000; // x = -30.4062, f(x) = 0.0000
    12'h867: soft_out = 32'h00000000; // x = -30.3906, f(x) = 0.0000
    12'h868: soft_out = 32'h00000000; // x = -30.3750, f(x) = 0.0000
    12'h869: soft_out = 32'h00000000; // x = -30.3594, f(x) = 0.0000
    12'h86A: soft_out = 32'h00000000; // x = -30.3438, f(x) = 0.0000
    12'h86B: soft_out = 32'h00000000; // x = -30.3281, f(x) = 0.0000
    12'h86C: soft_out = 32'h00000000; // x = -30.3125, f(x) = 0.0000
    12'h86D: soft_out = 32'h00000000; // x = -30.2969, f(x) = 0.0000
    12'h86E: soft_out = 32'h00000000; // x = -30.2812, f(x) = 0.0000
    12'h86F: soft_out = 32'h00000000; // x = -30.2656, f(x) = 0.0000
    12'h870: soft_out = 32'h00000000; // x = -30.2500, f(x) = 0.0000
    12'h871: soft_out = 32'h00000000; // x = -30.2344, f(x) = 0.0000
    12'h872: soft_out = 32'h00000000; // x = -30.2188, f(x) = 0.0000
    12'h873: soft_out = 32'h00000000; // x = -30.2031, f(x) = 0.0000
    12'h874: soft_out = 32'h00000000; // x = -30.1875, f(x) = 0.0000
    12'h875: soft_out = 32'h00000000; // x = -30.1719, f(x) = 0.0000
    12'h876: soft_out = 32'h00000000; // x = -30.1562, f(x) = 0.0000
    12'h877: soft_out = 32'h00000000; // x = -30.1406, f(x) = 0.0000
    12'h878: soft_out = 32'h00000000; // x = -30.1250, f(x) = 0.0000
    12'h879: soft_out = 32'h00000000; // x = -30.1094, f(x) = 0.0000
    12'h87A: soft_out = 32'h00000000; // x = -30.0938, f(x) = 0.0000
    12'h87B: soft_out = 32'h00000000; // x = -30.0781, f(x) = 0.0000
    12'h87C: soft_out = 32'h00000000; // x = -30.0625, f(x) = 0.0000
    12'h87D: soft_out = 32'h00000000; // x = -30.0469, f(x) = 0.0000
    12'h87E: soft_out = 32'h00000000; // x = -30.0312, f(x) = 0.0000
    12'h87F: soft_out = 32'h00000000; // x = -30.0156, f(x) = 0.0000
    12'h880: soft_out = 32'h00000000; // x = -30.0000, f(x) = 0.0000
    12'h881: soft_out = 32'h00000000; // x = -29.9844, f(x) = 0.0000
    12'h882: soft_out = 32'h00000000; // x = -29.9688, f(x) = 0.0000
    12'h883: soft_out = 32'h00000000; // x = -29.9531, f(x) = 0.0000
    12'h884: soft_out = 32'h00000000; // x = -29.9375, f(x) = 0.0000
    12'h885: soft_out = 32'h00000000; // x = -29.9219, f(x) = 0.0000
    12'h886: soft_out = 32'h00000000; // x = -29.9062, f(x) = 0.0000
    12'h887: soft_out = 32'h00000000; // x = -29.8906, f(x) = 0.0000
    12'h888: soft_out = 32'h00000000; // x = -29.8750, f(x) = 0.0000
    12'h889: soft_out = 32'h00000000; // x = -29.8594, f(x) = 0.0000
    12'h88A: soft_out = 32'h00000000; // x = -29.8438, f(x) = 0.0000
    12'h88B: soft_out = 32'h00000000; // x = -29.8281, f(x) = 0.0000
    12'h88C: soft_out = 32'h00000000; // x = -29.8125, f(x) = 0.0000
    12'h88D: soft_out = 32'h00000000; // x = -29.7969, f(x) = 0.0000
    12'h88E: soft_out = 32'h00000000; // x = -29.7812, f(x) = 0.0000
    12'h88F: soft_out = 32'h00000000; // x = -29.7656, f(x) = 0.0000
    12'h890: soft_out = 32'h00000000; // x = -29.7500, f(x) = 0.0000
    12'h891: soft_out = 32'h00000000; // x = -29.7344, f(x) = 0.0000
    12'h892: soft_out = 32'h00000000; // x = -29.7188, f(x) = 0.0000
    12'h893: soft_out = 32'h00000000; // x = -29.7031, f(x) = 0.0000
    12'h894: soft_out = 32'h00000000; // x = -29.6875, f(x) = 0.0000
    12'h895: soft_out = 32'h00000000; // x = -29.6719, f(x) = 0.0000
    12'h896: soft_out = 32'h00000000; // x = -29.6562, f(x) = 0.0000
    12'h897: soft_out = 32'h00000000; // x = -29.6406, f(x) = 0.0000
    12'h898: soft_out = 32'h00000000; // x = -29.6250, f(x) = 0.0000
    12'h899: soft_out = 32'h00000000; // x = -29.6094, f(x) = 0.0000
    12'h89A: soft_out = 32'h00000000; // x = -29.5938, f(x) = 0.0000
    12'h89B: soft_out = 32'h00000000; // x = -29.5781, f(x) = 0.0000
    12'h89C: soft_out = 32'h00000000; // x = -29.5625, f(x) = 0.0000
    12'h89D: soft_out = 32'h00000000; // x = -29.5469, f(x) = 0.0000
    12'h89E: soft_out = 32'h00000000; // x = -29.5312, f(x) = 0.0000
    12'h89F: soft_out = 32'h00000000; // x = -29.5156, f(x) = 0.0000
    12'h8A0: soft_out = 32'h00000000; // x = -29.5000, f(x) = 0.0000
    12'h8A1: soft_out = 32'h00000000; // x = -29.4844, f(x) = 0.0000
    12'h8A2: soft_out = 32'h00000000; // x = -29.4688, f(x) = 0.0000
    12'h8A3: soft_out = 32'h00000000; // x = -29.4531, f(x) = 0.0000
    12'h8A4: soft_out = 32'h00000000; // x = -29.4375, f(x) = 0.0000
    12'h8A5: soft_out = 32'h00000000; // x = -29.4219, f(x) = 0.0000
    12'h8A6: soft_out = 32'h00000000; // x = -29.4062, f(x) = 0.0000
    12'h8A7: soft_out = 32'h00000000; // x = -29.3906, f(x) = 0.0000
    12'h8A8: soft_out = 32'h00000000; // x = -29.3750, f(x) = 0.0000
    12'h8A9: soft_out = 32'h00000000; // x = -29.3594, f(x) = 0.0000
    12'h8AA: soft_out = 32'h00000000; // x = -29.3438, f(x) = 0.0000
    12'h8AB: soft_out = 32'h00000000; // x = -29.3281, f(x) = 0.0000
    12'h8AC: soft_out = 32'h00000000; // x = -29.3125, f(x) = 0.0000
    12'h8AD: soft_out = 32'h00000000; // x = -29.2969, f(x) = 0.0000
    12'h8AE: soft_out = 32'h00000000; // x = -29.2812, f(x) = 0.0000
    12'h8AF: soft_out = 32'h00000000; // x = -29.2656, f(x) = 0.0000
    12'h8B0: soft_out = 32'h00000000; // x = -29.2500, f(x) = 0.0000
    12'h8B1: soft_out = 32'h00000000; // x = -29.2344, f(x) = 0.0000
    12'h8B2: soft_out = 32'h00000000; // x = -29.2188, f(x) = 0.0000
    12'h8B3: soft_out = 32'h00000000; // x = -29.2031, f(x) = 0.0000
    12'h8B4: soft_out = 32'h00000000; // x = -29.1875, f(x) = 0.0000
    12'h8B5: soft_out = 32'h00000000; // x = -29.1719, f(x) = 0.0000
    12'h8B6: soft_out = 32'h00000000; // x = -29.1562, f(x) = 0.0000
    12'h8B7: soft_out = 32'h00000000; // x = -29.1406, f(x) = 0.0000
    12'h8B8: soft_out = 32'h00000000; // x = -29.1250, f(x) = 0.0000
    12'h8B9: soft_out = 32'h00000000; // x = -29.1094, f(x) = 0.0000
    12'h8BA: soft_out = 32'h00000000; // x = -29.0938, f(x) = 0.0000
    12'h8BB: soft_out = 32'h00000000; // x = -29.0781, f(x) = 0.0000
    12'h8BC: soft_out = 32'h00000000; // x = -29.0625, f(x) = 0.0000
    12'h8BD: soft_out = 32'h00000000; // x = -29.0469, f(x) = 0.0000
    12'h8BE: soft_out = 32'h00000000; // x = -29.0312, f(x) = 0.0000
    12'h8BF: soft_out = 32'h00000000; // x = -29.0156, f(x) = 0.0000
    12'h8C0: soft_out = 32'h00000000; // x = -29.0000, f(x) = 0.0000
    12'h8C1: soft_out = 32'h00000000; // x = -28.9844, f(x) = 0.0000
    12'h8C2: soft_out = 32'h00000000; // x = -28.9688, f(x) = 0.0000
    12'h8C3: soft_out = 32'h00000000; // x = -28.9531, f(x) = 0.0000
    12'h8C4: soft_out = 32'h00000000; // x = -28.9375, f(x) = 0.0000
    12'h8C5: soft_out = 32'h00000000; // x = -28.9219, f(x) = 0.0000
    12'h8C6: soft_out = 32'h00000000; // x = -28.9062, f(x) = 0.0000
    12'h8C7: soft_out = 32'h00000000; // x = -28.8906, f(x) = 0.0000
    12'h8C8: soft_out = 32'h00000000; // x = -28.8750, f(x) = 0.0000
    12'h8C9: soft_out = 32'h00000000; // x = -28.8594, f(x) = 0.0000
    12'h8CA: soft_out = 32'h00000000; // x = -28.8438, f(x) = 0.0000
    12'h8CB: soft_out = 32'h00000000; // x = -28.8281, f(x) = 0.0000
    12'h8CC: soft_out = 32'h00000000; // x = -28.8125, f(x) = 0.0000
    12'h8CD: soft_out = 32'h00000000; // x = -28.7969, f(x) = 0.0000
    12'h8CE: soft_out = 32'h00000000; // x = -28.7812, f(x) = 0.0000
    12'h8CF: soft_out = 32'h00000000; // x = -28.7656, f(x) = 0.0000
    12'h8D0: soft_out = 32'h00000000; // x = -28.7500, f(x) = 0.0000
    12'h8D1: soft_out = 32'h00000000; // x = -28.7344, f(x) = 0.0000
    12'h8D2: soft_out = 32'h00000000; // x = -28.7188, f(x) = 0.0000
    12'h8D3: soft_out = 32'h00000000; // x = -28.7031, f(x) = 0.0000
    12'h8D4: soft_out = 32'h00000000; // x = -28.6875, f(x) = 0.0000
    12'h8D5: soft_out = 32'h00000000; // x = -28.6719, f(x) = 0.0000
    12'h8D6: soft_out = 32'h00000000; // x = -28.6562, f(x) = 0.0000
    12'h8D7: soft_out = 32'h00000000; // x = -28.6406, f(x) = 0.0000
    12'h8D8: soft_out = 32'h00000000; // x = -28.6250, f(x) = 0.0000
    12'h8D9: soft_out = 32'h00000000; // x = -28.6094, f(x) = 0.0000
    12'h8DA: soft_out = 32'h00000000; // x = -28.5938, f(x) = 0.0000
    12'h8DB: soft_out = 32'h00000000; // x = -28.5781, f(x) = 0.0000
    12'h8DC: soft_out = 32'h00000000; // x = -28.5625, f(x) = 0.0000
    12'h8DD: soft_out = 32'h00000000; // x = -28.5469, f(x) = 0.0000
    12'h8DE: soft_out = 32'h00000000; // x = -28.5312, f(x) = 0.0000
    12'h8DF: soft_out = 32'h00000000; // x = -28.5156, f(x) = 0.0000
    12'h8E0: soft_out = 32'h00000000; // x = -28.5000, f(x) = 0.0000
    12'h8E1: soft_out = 32'h00000000; // x = -28.4844, f(x) = 0.0000
    12'h8E2: soft_out = 32'h00000000; // x = -28.4688, f(x) = 0.0000
    12'h8E3: soft_out = 32'h00000000; // x = -28.4531, f(x) = 0.0000
    12'h8E4: soft_out = 32'h00000000; // x = -28.4375, f(x) = 0.0000
    12'h8E5: soft_out = 32'h00000000; // x = -28.4219, f(x) = 0.0000
    12'h8E6: soft_out = 32'h00000000; // x = -28.4062, f(x) = 0.0000
    12'h8E7: soft_out = 32'h00000000; // x = -28.3906, f(x) = 0.0000
    12'h8E8: soft_out = 32'h00000000; // x = -28.3750, f(x) = 0.0000
    12'h8E9: soft_out = 32'h00000000; // x = -28.3594, f(x) = 0.0000
    12'h8EA: soft_out = 32'h00000000; // x = -28.3438, f(x) = 0.0000
    12'h8EB: soft_out = 32'h00000000; // x = -28.3281, f(x) = 0.0000
    12'h8EC: soft_out = 32'h00000000; // x = -28.3125, f(x) = 0.0000
    12'h8ED: soft_out = 32'h00000000; // x = -28.2969, f(x) = 0.0000
    12'h8EE: soft_out = 32'h00000000; // x = -28.2812, f(x) = 0.0000
    12'h8EF: soft_out = 32'h00000000; // x = -28.2656, f(x) = 0.0000
    12'h8F0: soft_out = 32'h00000000; // x = -28.2500, f(x) = 0.0000
    12'h8F1: soft_out = 32'h00000000; // x = -28.2344, f(x) = 0.0000
    12'h8F2: soft_out = 32'h00000000; // x = -28.2188, f(x) = 0.0000
    12'h8F3: soft_out = 32'h00000000; // x = -28.2031, f(x) = 0.0000
    12'h8F4: soft_out = 32'h00000000; // x = -28.1875, f(x) = 0.0000
    12'h8F5: soft_out = 32'h00000000; // x = -28.1719, f(x) = 0.0000
    12'h8F6: soft_out = 32'h00000000; // x = -28.1562, f(x) = 0.0000
    12'h8F7: soft_out = 32'h00000000; // x = -28.1406, f(x) = 0.0000
    12'h8F8: soft_out = 32'h00000000; // x = -28.1250, f(x) = 0.0000
    12'h8F9: soft_out = 32'h00000000; // x = -28.1094, f(x) = 0.0000
    12'h8FA: soft_out = 32'h00000000; // x = -28.0938, f(x) = 0.0000
    12'h8FB: soft_out = 32'h00000000; // x = -28.0781, f(x) = 0.0000
    12'h8FC: soft_out = 32'h00000000; // x = -28.0625, f(x) = 0.0000
    12'h8FD: soft_out = 32'h00000000; // x = -28.0469, f(x) = 0.0000
    12'h8FE: soft_out = 32'h00000000; // x = -28.0312, f(x) = 0.0000
    12'h8FF: soft_out = 32'h00000000; // x = -28.0156, f(x) = 0.0000
    12'h900: soft_out = 32'h00000000; // x = -28.0000, f(x) = 0.0000
    12'h901: soft_out = 32'h00000000; // x = -27.9844, f(x) = 0.0000
    12'h902: soft_out = 32'h00000000; // x = -27.9688, f(x) = 0.0000
    12'h903: soft_out = 32'h00000000; // x = -27.9531, f(x) = 0.0000
    12'h904: soft_out = 32'h00000000; // x = -27.9375, f(x) = 0.0000
    12'h905: soft_out = 32'h00000000; // x = -27.9219, f(x) = 0.0000
    12'h906: soft_out = 32'h00000000; // x = -27.9062, f(x) = 0.0000
    12'h907: soft_out = 32'h00000000; // x = -27.8906, f(x) = 0.0000
    12'h908: soft_out = 32'h00000000; // x = -27.8750, f(x) = 0.0000
    12'h909: soft_out = 32'h00000000; // x = -27.8594, f(x) = 0.0000
    12'h90A: soft_out = 32'h00000000; // x = -27.8438, f(x) = 0.0000
    12'h90B: soft_out = 32'h00000000; // x = -27.8281, f(x) = 0.0000
    12'h90C: soft_out = 32'h00000000; // x = -27.8125, f(x) = 0.0000
    12'h90D: soft_out = 32'h00000000; // x = -27.7969, f(x) = 0.0000
    12'h90E: soft_out = 32'h00000000; // x = -27.7812, f(x) = 0.0000
    12'h90F: soft_out = 32'h00000000; // x = -27.7656, f(x) = 0.0000
    12'h910: soft_out = 32'h00000000; // x = -27.7500, f(x) = 0.0000
    12'h911: soft_out = 32'h00000000; // x = -27.7344, f(x) = 0.0000
    12'h912: soft_out = 32'h00000000; // x = -27.7188, f(x) = 0.0000
    12'h913: soft_out = 32'h00000000; // x = -27.7031, f(x) = 0.0000
    12'h914: soft_out = 32'h00000000; // x = -27.6875, f(x) = 0.0000
    12'h915: soft_out = 32'h00000000; // x = -27.6719, f(x) = 0.0000
    12'h916: soft_out = 32'h00000000; // x = -27.6562, f(x) = 0.0000
    12'h917: soft_out = 32'h00000000; // x = -27.6406, f(x) = 0.0000
    12'h918: soft_out = 32'h00000000; // x = -27.6250, f(x) = 0.0000
    12'h919: soft_out = 32'h00000000; // x = -27.6094, f(x) = 0.0000
    12'h91A: soft_out = 32'h00000000; // x = -27.5938, f(x) = 0.0000
    12'h91B: soft_out = 32'h00000000; // x = -27.5781, f(x) = 0.0000
    12'h91C: soft_out = 32'h00000000; // x = -27.5625, f(x) = 0.0000
    12'h91D: soft_out = 32'h00000000; // x = -27.5469, f(x) = 0.0000
    12'h91E: soft_out = 32'h00000000; // x = -27.5312, f(x) = 0.0000
    12'h91F: soft_out = 32'h00000000; // x = -27.5156, f(x) = 0.0000
    12'h920: soft_out = 32'h00000000; // x = -27.5000, f(x) = 0.0000
    12'h921: soft_out = 32'h00000000; // x = -27.4844, f(x) = 0.0000
    12'h922: soft_out = 32'h00000000; // x = -27.4688, f(x) = 0.0000
    12'h923: soft_out = 32'h00000000; // x = -27.4531, f(x) = 0.0000
    12'h924: soft_out = 32'h00000000; // x = -27.4375, f(x) = 0.0000
    12'h925: soft_out = 32'h00000000; // x = -27.4219, f(x) = 0.0000
    12'h926: soft_out = 32'h00000000; // x = -27.4062, f(x) = 0.0000
    12'h927: soft_out = 32'h00000000; // x = -27.3906, f(x) = 0.0000
    12'h928: soft_out = 32'h00000000; // x = -27.3750, f(x) = 0.0000
    12'h929: soft_out = 32'h00000000; // x = -27.3594, f(x) = 0.0000
    12'h92A: soft_out = 32'h00000000; // x = -27.3438, f(x) = 0.0000
    12'h92B: soft_out = 32'h00000000; // x = -27.3281, f(x) = 0.0000
    12'h92C: soft_out = 32'h00000000; // x = -27.3125, f(x) = 0.0000
    12'h92D: soft_out = 32'h00000000; // x = -27.2969, f(x) = 0.0000
    12'h92E: soft_out = 32'h00000000; // x = -27.2812, f(x) = 0.0000
    12'h92F: soft_out = 32'h00000000; // x = -27.2656, f(x) = 0.0000
    12'h930: soft_out = 32'h00000000; // x = -27.2500, f(x) = 0.0000
    12'h931: soft_out = 32'h00000000; // x = -27.2344, f(x) = 0.0000
    12'h932: soft_out = 32'h00000000; // x = -27.2188, f(x) = 0.0000
    12'h933: soft_out = 32'h00000000; // x = -27.2031, f(x) = 0.0000
    12'h934: soft_out = 32'h00000000; // x = -27.1875, f(x) = 0.0000
    12'h935: soft_out = 32'h00000000; // x = -27.1719, f(x) = 0.0000
    12'h936: soft_out = 32'h00000000; // x = -27.1562, f(x) = 0.0000
    12'h937: soft_out = 32'h00000000; // x = -27.1406, f(x) = 0.0000
    12'h938: soft_out = 32'h00000000; // x = -27.1250, f(x) = 0.0000
    12'h939: soft_out = 32'h00000000; // x = -27.1094, f(x) = 0.0000
    12'h93A: soft_out = 32'h00000000; // x = -27.0938, f(x) = 0.0000
    12'h93B: soft_out = 32'h00000000; // x = -27.0781, f(x) = 0.0000
    12'h93C: soft_out = 32'h00000000; // x = -27.0625, f(x) = 0.0000
    12'h93D: soft_out = 32'h00000000; // x = -27.0469, f(x) = 0.0000
    12'h93E: soft_out = 32'h00000000; // x = -27.0312, f(x) = 0.0000
    12'h93F: soft_out = 32'h00000000; // x = -27.0156, f(x) = 0.0000
    12'h940: soft_out = 32'h00000000; // x = -27.0000, f(x) = 0.0000
    12'h941: soft_out = 32'h00000000; // x = -26.9844, f(x) = 0.0000
    12'h942: soft_out = 32'h00000000; // x = -26.9688, f(x) = 0.0000
    12'h943: soft_out = 32'h00000000; // x = -26.9531, f(x) = 0.0000
    12'h944: soft_out = 32'h00000000; // x = -26.9375, f(x) = 0.0000
    12'h945: soft_out = 32'h00000000; // x = -26.9219, f(x) = 0.0000
    12'h946: soft_out = 32'h00000000; // x = -26.9062, f(x) = 0.0000
    12'h947: soft_out = 32'h00000000; // x = -26.8906, f(x) = 0.0000
    12'h948: soft_out = 32'h00000000; // x = -26.8750, f(x) = 0.0000
    12'h949: soft_out = 32'h00000000; // x = -26.8594, f(x) = 0.0000
    12'h94A: soft_out = 32'h00000000; // x = -26.8438, f(x) = 0.0000
    12'h94B: soft_out = 32'h00000000; // x = -26.8281, f(x) = 0.0000
    12'h94C: soft_out = 32'h00000000; // x = -26.8125, f(x) = 0.0000
    12'h94D: soft_out = 32'h00000000; // x = -26.7969, f(x) = 0.0000
    12'h94E: soft_out = 32'h00000000; // x = -26.7812, f(x) = 0.0000
    12'h94F: soft_out = 32'h00000000; // x = -26.7656, f(x) = 0.0000
    12'h950: soft_out = 32'h00000000; // x = -26.7500, f(x) = 0.0000
    12'h951: soft_out = 32'h00000000; // x = -26.7344, f(x) = 0.0000
    12'h952: soft_out = 32'h00000000; // x = -26.7188, f(x) = 0.0000
    12'h953: soft_out = 32'h00000000; // x = -26.7031, f(x) = 0.0000
    12'h954: soft_out = 32'h00000000; // x = -26.6875, f(x) = 0.0000
    12'h955: soft_out = 32'h00000000; // x = -26.6719, f(x) = 0.0000
    12'h956: soft_out = 32'h00000000; // x = -26.6562, f(x) = 0.0000
    12'h957: soft_out = 32'h00000000; // x = -26.6406, f(x) = 0.0000
    12'h958: soft_out = 32'h00000000; // x = -26.6250, f(x) = 0.0000
    12'h959: soft_out = 32'h00000000; // x = -26.6094, f(x) = 0.0000
    12'h95A: soft_out = 32'h00000000; // x = -26.5938, f(x) = 0.0000
    12'h95B: soft_out = 32'h00000000; // x = -26.5781, f(x) = 0.0000
    12'h95C: soft_out = 32'h00000000; // x = -26.5625, f(x) = 0.0000
    12'h95D: soft_out = 32'h00000000; // x = -26.5469, f(x) = 0.0000
    12'h95E: soft_out = 32'h00000000; // x = -26.5312, f(x) = 0.0000
    12'h95F: soft_out = 32'h00000000; // x = -26.5156, f(x) = 0.0000
    12'h960: soft_out = 32'h00000000; // x = -26.5000, f(x) = 0.0000
    12'h961: soft_out = 32'h00000000; // x = -26.4844, f(x) = 0.0000
    12'h962: soft_out = 32'h00000000; // x = -26.4688, f(x) = 0.0000
    12'h963: soft_out = 32'h00000000; // x = -26.4531, f(x) = 0.0000
    12'h964: soft_out = 32'h00000000; // x = -26.4375, f(x) = 0.0000
    12'h965: soft_out = 32'h00000000; // x = -26.4219, f(x) = 0.0000
    12'h966: soft_out = 32'h00000000; // x = -26.4062, f(x) = 0.0000
    12'h967: soft_out = 32'h00000000; // x = -26.3906, f(x) = 0.0000
    12'h968: soft_out = 32'h00000000; // x = -26.3750, f(x) = 0.0000
    12'h969: soft_out = 32'h00000000; // x = -26.3594, f(x) = 0.0000
    12'h96A: soft_out = 32'h00000000; // x = -26.3438, f(x) = 0.0000
    12'h96B: soft_out = 32'h00000000; // x = -26.3281, f(x) = 0.0000
    12'h96C: soft_out = 32'h00000000; // x = -26.3125, f(x) = 0.0000
    12'h96D: soft_out = 32'h00000000; // x = -26.2969, f(x) = 0.0000
    12'h96E: soft_out = 32'h00000000; // x = -26.2812, f(x) = 0.0000
    12'h96F: soft_out = 32'h00000000; // x = -26.2656, f(x) = 0.0000
    12'h970: soft_out = 32'h00000000; // x = -26.2500, f(x) = 0.0000
    12'h971: soft_out = 32'h00000000; // x = -26.2344, f(x) = 0.0000
    12'h972: soft_out = 32'h00000000; // x = -26.2188, f(x) = 0.0000
    12'h973: soft_out = 32'h00000000; // x = -26.2031, f(x) = 0.0000
    12'h974: soft_out = 32'h00000000; // x = -26.1875, f(x) = 0.0000
    12'h975: soft_out = 32'h00000000; // x = -26.1719, f(x) = 0.0000
    12'h976: soft_out = 32'h00000000; // x = -26.1562, f(x) = 0.0000
    12'h977: soft_out = 32'h00000000; // x = -26.1406, f(x) = 0.0000
    12'h978: soft_out = 32'h00000000; // x = -26.1250, f(x) = 0.0000
    12'h979: soft_out = 32'h00000000; // x = -26.1094, f(x) = 0.0000
    12'h97A: soft_out = 32'h00000000; // x = -26.0938, f(x) = 0.0000
    12'h97B: soft_out = 32'h00000000; // x = -26.0781, f(x) = 0.0000
    12'h97C: soft_out = 32'h00000000; // x = -26.0625, f(x) = 0.0000
    12'h97D: soft_out = 32'h00000000; // x = -26.0469, f(x) = 0.0000
    12'h97E: soft_out = 32'h00000000; // x = -26.0312, f(x) = 0.0000
    12'h97F: soft_out = 32'h00000000; // x = -26.0156, f(x) = 0.0000
    12'h980: soft_out = 32'h00000000; // x = -26.0000, f(x) = 0.0000
    12'h981: soft_out = 32'h00000000; // x = -25.9844, f(x) = 0.0000
    12'h982: soft_out = 32'h00000000; // x = -25.9688, f(x) = 0.0000
    12'h983: soft_out = 32'h00000000; // x = -25.9531, f(x) = 0.0000
    12'h984: soft_out = 32'h00000000; // x = -25.9375, f(x) = 0.0000
    12'h985: soft_out = 32'h00000000; // x = -25.9219, f(x) = 0.0000
    12'h986: soft_out = 32'h00000000; // x = -25.9062, f(x) = 0.0000
    12'h987: soft_out = 32'h00000000; // x = -25.8906, f(x) = 0.0000
    12'h988: soft_out = 32'h00000000; // x = -25.8750, f(x) = 0.0000
    12'h989: soft_out = 32'h00000000; // x = -25.8594, f(x) = 0.0000
    12'h98A: soft_out = 32'h00000000; // x = -25.8438, f(x) = 0.0000
    12'h98B: soft_out = 32'h00000000; // x = -25.8281, f(x) = 0.0000
    12'h98C: soft_out = 32'h00000000; // x = -25.8125, f(x) = 0.0000
    12'h98D: soft_out = 32'h00000000; // x = -25.7969, f(x) = 0.0000
    12'h98E: soft_out = 32'h00000000; // x = -25.7812, f(x) = 0.0000
    12'h98F: soft_out = 32'h00000000; // x = -25.7656, f(x) = 0.0000
    12'h990: soft_out = 32'h00000000; // x = -25.7500, f(x) = 0.0000
    12'h991: soft_out = 32'h00000000; // x = -25.7344, f(x) = 0.0000
    12'h992: soft_out = 32'h00000000; // x = -25.7188, f(x) = 0.0000
    12'h993: soft_out = 32'h00000000; // x = -25.7031, f(x) = 0.0000
    12'h994: soft_out = 32'h00000000; // x = -25.6875, f(x) = 0.0000
    12'h995: soft_out = 32'h00000000; // x = -25.6719, f(x) = 0.0000
    12'h996: soft_out = 32'h00000000; // x = -25.6562, f(x) = 0.0000
    12'h997: soft_out = 32'h00000000; // x = -25.6406, f(x) = 0.0000
    12'h998: soft_out = 32'h00000000; // x = -25.6250, f(x) = 0.0000
    12'h999: soft_out = 32'h00000000; // x = -25.6094, f(x) = 0.0000
    12'h99A: soft_out = 32'h00000000; // x = -25.5938, f(x) = 0.0000
    12'h99B: soft_out = 32'h00000000; // x = -25.5781, f(x) = 0.0000
    12'h99C: soft_out = 32'h00000000; // x = -25.5625, f(x) = 0.0000
    12'h99D: soft_out = 32'h00000000; // x = -25.5469, f(x) = 0.0000
    12'h99E: soft_out = 32'h00000000; // x = -25.5312, f(x) = 0.0000
    12'h99F: soft_out = 32'h00000000; // x = -25.5156, f(x) = 0.0000
    12'h9A0: soft_out = 32'h00000000; // x = -25.5000, f(x) = 0.0000
    12'h9A1: soft_out = 32'h00000000; // x = -25.4844, f(x) = 0.0000
    12'h9A2: soft_out = 32'h00000000; // x = -25.4688, f(x) = 0.0000
    12'h9A3: soft_out = 32'h00000000; // x = -25.4531, f(x) = 0.0000
    12'h9A4: soft_out = 32'h00000000; // x = -25.4375, f(x) = 0.0000
    12'h9A5: soft_out = 32'h00000000; // x = -25.4219, f(x) = 0.0000
    12'h9A6: soft_out = 32'h00000000; // x = -25.4062, f(x) = 0.0000
    12'h9A7: soft_out = 32'h00000000; // x = -25.3906, f(x) = 0.0000
    12'h9A8: soft_out = 32'h00000000; // x = -25.3750, f(x) = 0.0000
    12'h9A9: soft_out = 32'h00000000; // x = -25.3594, f(x) = 0.0000
    12'h9AA: soft_out = 32'h00000000; // x = -25.3438, f(x) = 0.0000
    12'h9AB: soft_out = 32'h00000000; // x = -25.3281, f(x) = 0.0000
    12'h9AC: soft_out = 32'h00000000; // x = -25.3125, f(x) = 0.0000
    12'h9AD: soft_out = 32'h00000000; // x = -25.2969, f(x) = 0.0000
    12'h9AE: soft_out = 32'h00000000; // x = -25.2812, f(x) = 0.0000
    12'h9AF: soft_out = 32'h00000000; // x = -25.2656, f(x) = 0.0000
    12'h9B0: soft_out = 32'h00000000; // x = -25.2500, f(x) = 0.0000
    12'h9B1: soft_out = 32'h00000000; // x = -25.2344, f(x) = 0.0000
    12'h9B2: soft_out = 32'h00000000; // x = -25.2188, f(x) = 0.0000
    12'h9B3: soft_out = 32'h00000000; // x = -25.2031, f(x) = 0.0000
    12'h9B4: soft_out = 32'h00000000; // x = -25.1875, f(x) = 0.0000
    12'h9B5: soft_out = 32'h00000000; // x = -25.1719, f(x) = 0.0000
    12'h9B6: soft_out = 32'h00000000; // x = -25.1562, f(x) = 0.0000
    12'h9B7: soft_out = 32'h00000000; // x = -25.1406, f(x) = 0.0000
    12'h9B8: soft_out = 32'h00000000; // x = -25.1250, f(x) = 0.0000
    12'h9B9: soft_out = 32'h00000000; // x = -25.1094, f(x) = 0.0000
    12'h9BA: soft_out = 32'h00000000; // x = -25.0938, f(x) = 0.0000
    12'h9BB: soft_out = 32'h00000000; // x = -25.0781, f(x) = 0.0000
    12'h9BC: soft_out = 32'h00000000; // x = -25.0625, f(x) = 0.0000
    12'h9BD: soft_out = 32'h00000000; // x = -25.0469, f(x) = 0.0000
    12'h9BE: soft_out = 32'h00000000; // x = -25.0312, f(x) = 0.0000
    12'h9BF: soft_out = 32'h00000000; // x = -25.0156, f(x) = 0.0000
    12'h9C0: soft_out = 32'h00000000; // x = -25.0000, f(x) = 0.0000
    12'h9C1: soft_out = 32'h00000000; // x = -24.9844, f(x) = 0.0000
    12'h9C2: soft_out = 32'h00000000; // x = -24.9688, f(x) = 0.0000
    12'h9C3: soft_out = 32'h00000000; // x = -24.9531, f(x) = 0.0000
    12'h9C4: soft_out = 32'h00000000; // x = -24.9375, f(x) = 0.0000
    12'h9C5: soft_out = 32'h00000000; // x = -24.9219, f(x) = 0.0000
    12'h9C6: soft_out = 32'h00000000; // x = -24.9062, f(x) = 0.0000
    12'h9C7: soft_out = 32'h00000000; // x = -24.8906, f(x) = 0.0000
    12'h9C8: soft_out = 32'h00000000; // x = -24.8750, f(x) = 0.0000
    12'h9C9: soft_out = 32'h00000000; // x = -24.8594, f(x) = 0.0000
    12'h9CA: soft_out = 32'h00000000; // x = -24.8438, f(x) = 0.0000
    12'h9CB: soft_out = 32'h00000000; // x = -24.8281, f(x) = 0.0000
    12'h9CC: soft_out = 32'h00000000; // x = -24.8125, f(x) = 0.0000
    12'h9CD: soft_out = 32'h00000000; // x = -24.7969, f(x) = 0.0000
    12'h9CE: soft_out = 32'h00000000; // x = -24.7812, f(x) = 0.0000
    12'h9CF: soft_out = 32'h00000000; // x = -24.7656, f(x) = 0.0000
    12'h9D0: soft_out = 32'h00000000; // x = -24.7500, f(x) = 0.0000
    12'h9D1: soft_out = 32'h00000000; // x = -24.7344, f(x) = 0.0000
    12'h9D2: soft_out = 32'h00000000; // x = -24.7188, f(x) = 0.0000
    12'h9D3: soft_out = 32'h00000000; // x = -24.7031, f(x) = 0.0000
    12'h9D4: soft_out = 32'h00000000; // x = -24.6875, f(x) = 0.0000
    12'h9D5: soft_out = 32'h00000000; // x = -24.6719, f(x) = 0.0000
    12'h9D6: soft_out = 32'h00000000; // x = -24.6562, f(x) = 0.0000
    12'h9D7: soft_out = 32'h00000000; // x = -24.6406, f(x) = 0.0000
    12'h9D8: soft_out = 32'h00000000; // x = -24.6250, f(x) = 0.0000
    12'h9D9: soft_out = 32'h00000000; // x = -24.6094, f(x) = 0.0000
    12'h9DA: soft_out = 32'h00000000; // x = -24.5938, f(x) = 0.0000
    12'h9DB: soft_out = 32'h00000000; // x = -24.5781, f(x) = 0.0000
    12'h9DC: soft_out = 32'h00000000; // x = -24.5625, f(x) = 0.0000
    12'h9DD: soft_out = 32'h00000000; // x = -24.5469, f(x) = 0.0000
    12'h9DE: soft_out = 32'h00000000; // x = -24.5312, f(x) = 0.0000
    12'h9DF: soft_out = 32'h00000000; // x = -24.5156, f(x) = 0.0000
    12'h9E0: soft_out = 32'h00000000; // x = -24.5000, f(x) = 0.0000
    12'h9E1: soft_out = 32'h00000000; // x = -24.4844, f(x) = 0.0000
    12'h9E2: soft_out = 32'h00000000; // x = -24.4688, f(x) = 0.0000
    12'h9E3: soft_out = 32'h00000000; // x = -24.4531, f(x) = 0.0000
    12'h9E4: soft_out = 32'h00000000; // x = -24.4375, f(x) = 0.0000
    12'h9E5: soft_out = 32'h00000000; // x = -24.4219, f(x) = 0.0000
    12'h9E6: soft_out = 32'h00000000; // x = -24.4062, f(x) = 0.0000
    12'h9E7: soft_out = 32'h00000000; // x = -24.3906, f(x) = 0.0000
    12'h9E8: soft_out = 32'h00000000; // x = -24.3750, f(x) = 0.0000
    12'h9E9: soft_out = 32'h00000000; // x = -24.3594, f(x) = 0.0000
    12'h9EA: soft_out = 32'h00000000; // x = -24.3438, f(x) = 0.0000
    12'h9EB: soft_out = 32'h00000000; // x = -24.3281, f(x) = 0.0000
    12'h9EC: soft_out = 32'h00000000; // x = -24.3125, f(x) = 0.0000
    12'h9ED: soft_out = 32'h00000000; // x = -24.2969, f(x) = 0.0000
    12'h9EE: soft_out = 32'h00000000; // x = -24.2812, f(x) = 0.0000
    12'h9EF: soft_out = 32'h00000000; // x = -24.2656, f(x) = 0.0000
    12'h9F0: soft_out = 32'h00000000; // x = -24.2500, f(x) = 0.0000
    12'h9F1: soft_out = 32'h00000000; // x = -24.2344, f(x) = 0.0000
    12'h9F2: soft_out = 32'h00000000; // x = -24.2188, f(x) = 0.0000
    12'h9F3: soft_out = 32'h00000000; // x = -24.2031, f(x) = 0.0000
    12'h9F4: soft_out = 32'h00000000; // x = -24.1875, f(x) = 0.0000
    12'h9F5: soft_out = 32'h00000000; // x = -24.1719, f(x) = 0.0000
    12'h9F6: soft_out = 32'h00000000; // x = -24.1562, f(x) = 0.0000
    12'h9F7: soft_out = 32'h00000000; // x = -24.1406, f(x) = 0.0000
    12'h9F8: soft_out = 32'h00000000; // x = -24.1250, f(x) = 0.0000
    12'h9F9: soft_out = 32'h00000000; // x = -24.1094, f(x) = 0.0000
    12'h9FA: soft_out = 32'h00000000; // x = -24.0938, f(x) = 0.0000
    12'h9FB: soft_out = 32'h00000000; // x = -24.0781, f(x) = 0.0000
    12'h9FC: soft_out = 32'h00000000; // x = -24.0625, f(x) = 0.0000
    12'h9FD: soft_out = 32'h00000000; // x = -24.0469, f(x) = 0.0000
    12'h9FE: soft_out = 32'h00000000; // x = -24.0312, f(x) = 0.0000
    12'h9FF: soft_out = 32'h00000000; // x = -24.0156, f(x) = 0.0000
    12'hA00: soft_out = 32'h00000000; // x = -24.0000, f(x) = 0.0000
    12'hA01: soft_out = 32'h00000000; // x = -23.9844, f(x) = 0.0000
    12'hA02: soft_out = 32'h00000000; // x = -23.9688, f(x) = 0.0000
    12'hA03: soft_out = 32'h00000000; // x = -23.9531, f(x) = 0.0000
    12'hA04: soft_out = 32'h00000000; // x = -23.9375, f(x) = 0.0000
    12'hA05: soft_out = 32'h00000000; // x = -23.9219, f(x) = 0.0000
    12'hA06: soft_out = 32'h00000000; // x = -23.9062, f(x) = 0.0000
    12'hA07: soft_out = 32'h00000000; // x = -23.8906, f(x) = 0.0000
    12'hA08: soft_out = 32'h00000000; // x = -23.8750, f(x) = 0.0000
    12'hA09: soft_out = 32'h00000000; // x = -23.8594, f(x) = 0.0000
    12'hA0A: soft_out = 32'h00000000; // x = -23.8438, f(x) = 0.0000
    12'hA0B: soft_out = 32'h00000000; // x = -23.8281, f(x) = 0.0000
    12'hA0C: soft_out = 32'h00000000; // x = -23.8125, f(x) = 0.0000
    12'hA0D: soft_out = 32'h00000000; // x = -23.7969, f(x) = 0.0000
    12'hA0E: soft_out = 32'h00000000; // x = -23.7812, f(x) = 0.0000
    12'hA0F: soft_out = 32'h00000000; // x = -23.7656, f(x) = 0.0000
    12'hA10: soft_out = 32'h00000000; // x = -23.7500, f(x) = 0.0000
    12'hA11: soft_out = 32'h00000000; // x = -23.7344, f(x) = 0.0000
    12'hA12: soft_out = 32'h00000000; // x = -23.7188, f(x) = 0.0000
    12'hA13: soft_out = 32'h00000000; // x = -23.7031, f(x) = 0.0000
    12'hA14: soft_out = 32'h00000000; // x = -23.6875, f(x) = 0.0000
    12'hA15: soft_out = 32'h00000000; // x = -23.6719, f(x) = 0.0000
    12'hA16: soft_out = 32'h00000000; // x = -23.6562, f(x) = 0.0000
    12'hA17: soft_out = 32'h00000000; // x = -23.6406, f(x) = 0.0000
    12'hA18: soft_out = 32'h00000000; // x = -23.6250, f(x) = 0.0000
    12'hA19: soft_out = 32'h00000000; // x = -23.6094, f(x) = 0.0000
    12'hA1A: soft_out = 32'h00000000; // x = -23.5938, f(x) = 0.0000
    12'hA1B: soft_out = 32'h00000000; // x = -23.5781, f(x) = 0.0000
    12'hA1C: soft_out = 32'h00000000; // x = -23.5625, f(x) = 0.0000
    12'hA1D: soft_out = 32'h00000000; // x = -23.5469, f(x) = 0.0000
    12'hA1E: soft_out = 32'h00000000; // x = -23.5312, f(x) = 0.0000
    12'hA1F: soft_out = 32'h00000000; // x = -23.5156, f(x) = 0.0000
    12'hA20: soft_out = 32'h00000000; // x = -23.5000, f(x) = 0.0000
    12'hA21: soft_out = 32'h00000000; // x = -23.4844, f(x) = 0.0000
    12'hA22: soft_out = 32'h00000000; // x = -23.4688, f(x) = 0.0000
    12'hA23: soft_out = 32'h00000000; // x = -23.4531, f(x) = 0.0000
    12'hA24: soft_out = 32'h00000000; // x = -23.4375, f(x) = 0.0000
    12'hA25: soft_out = 32'h00000000; // x = -23.4219, f(x) = 0.0000
    12'hA26: soft_out = 32'h00000000; // x = -23.4062, f(x) = 0.0000
    12'hA27: soft_out = 32'h00000000; // x = -23.3906, f(x) = 0.0000
    12'hA28: soft_out = 32'h00000000; // x = -23.3750, f(x) = 0.0000
    12'hA29: soft_out = 32'h00000000; // x = -23.3594, f(x) = 0.0000
    12'hA2A: soft_out = 32'h00000000; // x = -23.3438, f(x) = 0.0000
    12'hA2B: soft_out = 32'h00000000; // x = -23.3281, f(x) = 0.0000
    12'hA2C: soft_out = 32'h00000000; // x = -23.3125, f(x) = 0.0000
    12'hA2D: soft_out = 32'h00000000; // x = -23.2969, f(x) = 0.0000
    12'hA2E: soft_out = 32'h00000000; // x = -23.2812, f(x) = 0.0000
    12'hA2F: soft_out = 32'h00000000; // x = -23.2656, f(x) = 0.0000
    12'hA30: soft_out = 32'h00000000; // x = -23.2500, f(x) = 0.0000
    12'hA31: soft_out = 32'h00000000; // x = -23.2344, f(x) = 0.0000
    12'hA32: soft_out = 32'h00000000; // x = -23.2188, f(x) = 0.0000
    12'hA33: soft_out = 32'h00000000; // x = -23.2031, f(x) = 0.0000
    12'hA34: soft_out = 32'h00000000; // x = -23.1875, f(x) = 0.0000
    12'hA35: soft_out = 32'h00000000; // x = -23.1719, f(x) = 0.0000
    12'hA36: soft_out = 32'h00000000; // x = -23.1562, f(x) = 0.0000
    12'hA37: soft_out = 32'h00000000; // x = -23.1406, f(x) = 0.0000
    12'hA38: soft_out = 32'h00000000; // x = -23.1250, f(x) = 0.0000
    12'hA39: soft_out = 32'h00000000; // x = -23.1094, f(x) = 0.0000
    12'hA3A: soft_out = 32'h00000000; // x = -23.0938, f(x) = 0.0000
    12'hA3B: soft_out = 32'h00000000; // x = -23.0781, f(x) = 0.0000
    12'hA3C: soft_out = 32'h00000000; // x = -23.0625, f(x) = 0.0000
    12'hA3D: soft_out = 32'h00000000; // x = -23.0469, f(x) = 0.0000
    12'hA3E: soft_out = 32'h00000000; // x = -23.0312, f(x) = 0.0000
    12'hA3F: soft_out = 32'h00000000; // x = -23.0156, f(x) = 0.0000
    12'hA40: soft_out = 32'h00000000; // x = -23.0000, f(x) = 0.0000
    12'hA41: soft_out = 32'h00000000; // x = -22.9844, f(x) = 0.0000
    12'hA42: soft_out = 32'h00000000; // x = -22.9688, f(x) = 0.0000
    12'hA43: soft_out = 32'h00000000; // x = -22.9531, f(x) = 0.0000
    12'hA44: soft_out = 32'h00000000; // x = -22.9375, f(x) = 0.0000
    12'hA45: soft_out = 32'h00000000; // x = -22.9219, f(x) = 0.0000
    12'hA46: soft_out = 32'h00000000; // x = -22.9062, f(x) = 0.0000
    12'hA47: soft_out = 32'h00000000; // x = -22.8906, f(x) = 0.0000
    12'hA48: soft_out = 32'h00000000; // x = -22.8750, f(x) = 0.0000
    12'hA49: soft_out = 32'h00000000; // x = -22.8594, f(x) = 0.0000
    12'hA4A: soft_out = 32'h00000000; // x = -22.8438, f(x) = 0.0000
    12'hA4B: soft_out = 32'h00000000; // x = -22.8281, f(x) = 0.0000
    12'hA4C: soft_out = 32'h00000000; // x = -22.8125, f(x) = 0.0000
    12'hA4D: soft_out = 32'h00000000; // x = -22.7969, f(x) = 0.0000
    12'hA4E: soft_out = 32'h00000000; // x = -22.7812, f(x) = 0.0000
    12'hA4F: soft_out = 32'h00000000; // x = -22.7656, f(x) = 0.0000
    12'hA50: soft_out = 32'h00000000; // x = -22.7500, f(x) = 0.0000
    12'hA51: soft_out = 32'h00000000; // x = -22.7344, f(x) = 0.0000
    12'hA52: soft_out = 32'h00000000; // x = -22.7188, f(x) = 0.0000
    12'hA53: soft_out = 32'h00000000; // x = -22.7031, f(x) = 0.0000
    12'hA54: soft_out = 32'h00000000; // x = -22.6875, f(x) = 0.0000
    12'hA55: soft_out = 32'h00000000; // x = -22.6719, f(x) = 0.0000
    12'hA56: soft_out = 32'h00000000; // x = -22.6562, f(x) = 0.0000
    12'hA57: soft_out = 32'h00000000; // x = -22.6406, f(x) = 0.0000
    12'hA58: soft_out = 32'h00000000; // x = -22.6250, f(x) = 0.0000
    12'hA59: soft_out = 32'h00000000; // x = -22.6094, f(x) = 0.0000
    12'hA5A: soft_out = 32'h00000000; // x = -22.5938, f(x) = 0.0000
    12'hA5B: soft_out = 32'h00000000; // x = -22.5781, f(x) = 0.0000
    12'hA5C: soft_out = 32'h00000000; // x = -22.5625, f(x) = 0.0000
    12'hA5D: soft_out = 32'h00000000; // x = -22.5469, f(x) = 0.0000
    12'hA5E: soft_out = 32'h00000000; // x = -22.5312, f(x) = 0.0000
    12'hA5F: soft_out = 32'h00000000; // x = -22.5156, f(x) = 0.0000
    12'hA60: soft_out = 32'h00000000; // x = -22.5000, f(x) = 0.0000
    12'hA61: soft_out = 32'h00000000; // x = -22.4844, f(x) = 0.0000
    12'hA62: soft_out = 32'h00000000; // x = -22.4688, f(x) = 0.0000
    12'hA63: soft_out = 32'h00000000; // x = -22.4531, f(x) = 0.0000
    12'hA64: soft_out = 32'h00000000; // x = -22.4375, f(x) = 0.0000
    12'hA65: soft_out = 32'h00000000; // x = -22.4219, f(x) = 0.0000
    12'hA66: soft_out = 32'h00000000; // x = -22.4062, f(x) = 0.0000
    12'hA67: soft_out = 32'h00000000; // x = -22.3906, f(x) = 0.0000
    12'hA68: soft_out = 32'h00000000; // x = -22.3750, f(x) = 0.0000
    12'hA69: soft_out = 32'h00000000; // x = -22.3594, f(x) = 0.0000
    12'hA6A: soft_out = 32'h00000000; // x = -22.3438, f(x) = 0.0000
    12'hA6B: soft_out = 32'h00000000; // x = -22.3281, f(x) = 0.0000
    12'hA6C: soft_out = 32'h00000000; // x = -22.3125, f(x) = 0.0000
    12'hA6D: soft_out = 32'h00000000; // x = -22.2969, f(x) = 0.0000
    12'hA6E: soft_out = 32'h00000000; // x = -22.2812, f(x) = 0.0000
    12'hA6F: soft_out = 32'h00000000; // x = -22.2656, f(x) = 0.0000
    12'hA70: soft_out = 32'h00000000; // x = -22.2500, f(x) = 0.0000
    12'hA71: soft_out = 32'h00000000; // x = -22.2344, f(x) = 0.0000
    12'hA72: soft_out = 32'h00000000; // x = -22.2188, f(x) = 0.0000
    12'hA73: soft_out = 32'h00000000; // x = -22.2031, f(x) = 0.0000
    12'hA74: soft_out = 32'h00000000; // x = -22.1875, f(x) = 0.0000
    12'hA75: soft_out = 32'h00000001; // x = -22.1719, f(x) = 0.0000
    12'hA76: soft_out = 32'h00000001; // x = -22.1562, f(x) = 0.0000
    12'hA77: soft_out = 32'h00000001; // x = -22.1406, f(x) = 0.0000
    12'hA78: soft_out = 32'h00000001; // x = -22.1250, f(x) = 0.0000
    12'hA79: soft_out = 32'h00000001; // x = -22.1094, f(x) = 0.0000
    12'hA7A: soft_out = 32'h00000001; // x = -22.0938, f(x) = 0.0000
    12'hA7B: soft_out = 32'h00000001; // x = -22.0781, f(x) = 0.0000
    12'hA7C: soft_out = 32'h00000001; // x = -22.0625, f(x) = 0.0000
    12'hA7D: soft_out = 32'h00000001; // x = -22.0469, f(x) = 0.0000
    12'hA7E: soft_out = 32'h00000001; // x = -22.0312, f(x) = 0.0000
    12'hA7F: soft_out = 32'h00000001; // x = -22.0156, f(x) = 0.0000
    12'hA80: soft_out = 32'h00000001; // x = -22.0000, f(x) = 0.0000
    12'hA81: soft_out = 32'h00000001; // x = -21.9844, f(x) = 0.0000
    12'hA82: soft_out = 32'h00000001; // x = -21.9688, f(x) = 0.0000
    12'hA83: soft_out = 32'h00000001; // x = -21.9531, f(x) = 0.0000
    12'hA84: soft_out = 32'h00000001; // x = -21.9375, f(x) = 0.0000
    12'hA85: soft_out = 32'h00000001; // x = -21.9219, f(x) = 0.0000
    12'hA86: soft_out = 32'h00000001; // x = -21.9062, f(x) = 0.0000
    12'hA87: soft_out = 32'h00000001; // x = -21.8906, f(x) = 0.0000
    12'hA88: soft_out = 32'h00000001; // x = -21.8750, f(x) = 0.0000
    12'hA89: soft_out = 32'h00000001; // x = -21.8594, f(x) = 0.0000
    12'hA8A: soft_out = 32'h00000001; // x = -21.8438, f(x) = 0.0000
    12'hA8B: soft_out = 32'h00000001; // x = -21.8281, f(x) = 0.0000
    12'hA8C: soft_out = 32'h00000001; // x = -21.8125, f(x) = 0.0000
    12'hA8D: soft_out = 32'h00000001; // x = -21.7969, f(x) = 0.0000
    12'hA8E: soft_out = 32'h00000001; // x = -21.7812, f(x) = 0.0000
    12'hA8F: soft_out = 32'h00000001; // x = -21.7656, f(x) = 0.0000
    12'hA90: soft_out = 32'h00000001; // x = -21.7500, f(x) = 0.0000
    12'hA91: soft_out = 32'h00000001; // x = -21.7344, f(x) = 0.0000
    12'hA92: soft_out = 32'h00000001; // x = -21.7188, f(x) = 0.0000
    12'hA93: soft_out = 32'h00000001; // x = -21.7031, f(x) = 0.0000
    12'hA94: soft_out = 32'h00000001; // x = -21.6875, f(x) = 0.0000
    12'hA95: soft_out = 32'h00000001; // x = -21.6719, f(x) = 0.0000
    12'hA96: soft_out = 32'h00000001; // x = -21.6562, f(x) = 0.0000
    12'hA97: soft_out = 32'h00000001; // x = -21.6406, f(x) = 0.0000
    12'hA98: soft_out = 32'h00000001; // x = -21.6250, f(x) = 0.0000
    12'hA99: soft_out = 32'h00000001; // x = -21.6094, f(x) = 0.0000
    12'hA9A: soft_out = 32'h00000001; // x = -21.5938, f(x) = 0.0000
    12'hA9B: soft_out = 32'h00000001; // x = -21.5781, f(x) = 0.0000
    12'hA9C: soft_out = 32'h00000001; // x = -21.5625, f(x) = 0.0000
    12'hA9D: soft_out = 32'h00000001; // x = -21.5469, f(x) = 0.0000
    12'hA9E: soft_out = 32'h00000001; // x = -21.5312, f(x) = 0.0000
    12'hA9F: soft_out = 32'h00000001; // x = -21.5156, f(x) = 0.0000
    12'hAA0: soft_out = 32'h00000001; // x = -21.5000, f(x) = 0.0000
    12'hAA1: soft_out = 32'h00000001; // x = -21.4844, f(x) = 0.0000
    12'hAA2: soft_out = 32'h00000001; // x = -21.4688, f(x) = 0.0000
    12'hAA3: soft_out = 32'h00000001; // x = -21.4531, f(x) = 0.0000
    12'hAA4: soft_out = 32'h00000001; // x = -21.4375, f(x) = 0.0000
    12'hAA5: soft_out = 32'h00000001; // x = -21.4219, f(x) = 0.0000
    12'hAA6: soft_out = 32'h00000001; // x = -21.4062, f(x) = 0.0000
    12'hAA7: soft_out = 32'h00000001; // x = -21.3906, f(x) = 0.0000
    12'hAA8: soft_out = 32'h00000001; // x = -21.3750, f(x) = 0.0000
    12'hAA9: soft_out = 32'h00000001; // x = -21.3594, f(x) = 0.0000
    12'hAAA: soft_out = 32'h00000001; // x = -21.3438, f(x) = 0.0000
    12'hAAB: soft_out = 32'h00000001; // x = -21.3281, f(x) = 0.0000
    12'hAAC: soft_out = 32'h00000001; // x = -21.3125, f(x) = 0.0000
    12'hAAD: soft_out = 32'h00000001; // x = -21.2969, f(x) = 0.0000
    12'hAAE: soft_out = 32'h00000001; // x = -21.2812, f(x) = 0.0000
    12'hAAF: soft_out = 32'h00000001; // x = -21.2656, f(x) = 0.0000
    12'hAB0: soft_out = 32'h00000001; // x = -21.2500, f(x) = 0.0000
    12'hAB1: soft_out = 32'h00000001; // x = -21.2344, f(x) = 0.0000
    12'hAB2: soft_out = 32'h00000001; // x = -21.2188, f(x) = 0.0000
    12'hAB3: soft_out = 32'h00000001; // x = -21.2031, f(x) = 0.0000
    12'hAB4: soft_out = 32'h00000001; // x = -21.1875, f(x) = 0.0000
    12'hAB5: soft_out = 32'h00000001; // x = -21.1719, f(x) = 0.0000
    12'hAB6: soft_out = 32'h00000001; // x = -21.1562, f(x) = 0.0000
    12'hAB7: soft_out = 32'h00000001; // x = -21.1406, f(x) = 0.0000
    12'hAB8: soft_out = 32'h00000001; // x = -21.1250, f(x) = 0.0000
    12'hAB9: soft_out = 32'h00000001; // x = -21.1094, f(x) = 0.0000
    12'hABA: soft_out = 32'h00000001; // x = -21.0938, f(x) = 0.0000
    12'hABB: soft_out = 32'h00000002; // x = -21.0781, f(x) = 0.0000
    12'hABC: soft_out = 32'h00000002; // x = -21.0625, f(x) = 0.0000
    12'hABD: soft_out = 32'h00000002; // x = -21.0469, f(x) = 0.0000
    12'hABE: soft_out = 32'h00000002; // x = -21.0312, f(x) = 0.0000
    12'hABF: soft_out = 32'h00000002; // x = -21.0156, f(x) = 0.0000
    12'hAC0: soft_out = 32'h00000002; // x = -21.0000, f(x) = 0.0000
    12'hAC1: soft_out = 32'h00000002; // x = -20.9844, f(x) = 0.0000
    12'hAC2: soft_out = 32'h00000002; // x = -20.9688, f(x) = 0.0000
    12'hAC3: soft_out = 32'h00000002; // x = -20.9531, f(x) = 0.0000
    12'hAC4: soft_out = 32'h00000002; // x = -20.9375, f(x) = 0.0000
    12'hAC5: soft_out = 32'h00000002; // x = -20.9219, f(x) = 0.0000
    12'hAC6: soft_out = 32'h00000002; // x = -20.9062, f(x) = 0.0000
    12'hAC7: soft_out = 32'h00000002; // x = -20.8906, f(x) = 0.0000
    12'hAC8: soft_out = 32'h00000002; // x = -20.8750, f(x) = 0.0000
    12'hAC9: soft_out = 32'h00000002; // x = -20.8594, f(x) = 0.0000
    12'hACA: soft_out = 32'h00000002; // x = -20.8438, f(x) = 0.0000
    12'hACB: soft_out = 32'h00000002; // x = -20.8281, f(x) = 0.0000
    12'hACC: soft_out = 32'h00000002; // x = -20.8125, f(x) = 0.0000
    12'hACD: soft_out = 32'h00000002; // x = -20.7969, f(x) = 0.0000
    12'hACE: soft_out = 32'h00000002; // x = -20.7812, f(x) = 0.0000
    12'hACF: soft_out = 32'h00000002; // x = -20.7656, f(x) = 0.0000
    12'hAD0: soft_out = 32'h00000002; // x = -20.7500, f(x) = 0.0000
    12'hAD1: soft_out = 32'h00000002; // x = -20.7344, f(x) = 0.0000
    12'hAD2: soft_out = 32'h00000002; // x = -20.7188, f(x) = 0.0000
    12'hAD3: soft_out = 32'h00000002; // x = -20.7031, f(x) = 0.0000
    12'hAD4: soft_out = 32'h00000002; // x = -20.6875, f(x) = 0.0000
    12'hAD5: soft_out = 32'h00000002; // x = -20.6719, f(x) = 0.0000
    12'hAD6: soft_out = 32'h00000002; // x = -20.6562, f(x) = 0.0000
    12'hAD7: soft_out = 32'h00000002; // x = -20.6406, f(x) = 0.0000
    12'hAD8: soft_out = 32'h00000002; // x = -20.6250, f(x) = 0.0000
    12'hAD9: soft_out = 32'h00000002; // x = -20.6094, f(x) = 0.0000
    12'hADA: soft_out = 32'h00000002; // x = -20.5938, f(x) = 0.0000
    12'hADB: soft_out = 32'h00000002; // x = -20.5781, f(x) = 0.0000
    12'hADC: soft_out = 32'h00000003; // x = -20.5625, f(x) = 0.0000
    12'hADD: soft_out = 32'h00000003; // x = -20.5469, f(x) = 0.0000
    12'hADE: soft_out = 32'h00000003; // x = -20.5312, f(x) = 0.0000
    12'hADF: soft_out = 32'h00000003; // x = -20.5156, f(x) = 0.0000
    12'hAE0: soft_out = 32'h00000003; // x = -20.5000, f(x) = 0.0000
    12'hAE1: soft_out = 32'h00000003; // x = -20.4844, f(x) = 0.0000
    12'hAE2: soft_out = 32'h00000003; // x = -20.4688, f(x) = 0.0000
    12'hAE3: soft_out = 32'h00000003; // x = -20.4531, f(x) = 0.0000
    12'hAE4: soft_out = 32'h00000003; // x = -20.4375, f(x) = 0.0000
    12'hAE5: soft_out = 32'h00000003; // x = -20.4219, f(x) = 0.0000
    12'hAE6: soft_out = 32'h00000003; // x = -20.4062, f(x) = 0.0000
    12'hAE7: soft_out = 32'h00000003; // x = -20.3906, f(x) = 0.0000
    12'hAE8: soft_out = 32'h00000003; // x = -20.3750, f(x) = 0.0000
    12'hAE9: soft_out = 32'h00000003; // x = -20.3594, f(x) = 0.0000
    12'hAEA: soft_out = 32'h00000003; // x = -20.3438, f(x) = 0.0000
    12'hAEB: soft_out = 32'h00000003; // x = -20.3281, f(x) = 0.0000
    12'hAEC: soft_out = 32'h00000003; // x = -20.3125, f(x) = 0.0000
    12'hAED: soft_out = 32'h00000003; // x = -20.2969, f(x) = 0.0000
    12'hAEE: soft_out = 32'h00000003; // x = -20.2812, f(x) = 0.0000
    12'hAEF: soft_out = 32'h00000003; // x = -20.2656, f(x) = 0.0000
    12'hAF0: soft_out = 32'h00000003; // x = -20.2500, f(x) = 0.0000
    12'hAF1: soft_out = 32'h00000004; // x = -20.2344, f(x) = 0.0000
    12'hAF2: soft_out = 32'h00000004; // x = -20.2188, f(x) = 0.0000
    12'hAF3: soft_out = 32'h00000004; // x = -20.2031, f(x) = 0.0000
    12'hAF4: soft_out = 32'h00000004; // x = -20.1875, f(x) = 0.0000
    12'hAF5: soft_out = 32'h00000004; // x = -20.1719, f(x) = 0.0000
    12'hAF6: soft_out = 32'h00000004; // x = -20.1562, f(x) = 0.0000
    12'hAF7: soft_out = 32'h00000004; // x = -20.1406, f(x) = 0.0000
    12'hAF8: soft_out = 32'h00000004; // x = -20.1250, f(x) = 0.0000
    12'hAF9: soft_out = 32'h00000004; // x = -20.1094, f(x) = 0.0000
    12'hAFA: soft_out = 32'h00000004; // x = -20.0938, f(x) = 0.0000
    12'hAFB: soft_out = 32'h00000004; // x = -20.0781, f(x) = 0.0000
    12'hAFC: soft_out = 32'h00000004; // x = -20.0625, f(x) = 0.0000
    12'hAFD: soft_out = 32'h00000004; // x = -20.0469, f(x) = 0.0000
    12'hAFE: soft_out = 32'h00000004; // x = -20.0312, f(x) = 0.0000
    12'hAFF: soft_out = 32'h00000004; // x = -20.0156, f(x) = 0.0000
    12'hB00: soft_out = 32'h00000004; // x = -20.0000, f(x) = 0.0000
    12'hB01: soft_out = 32'h00000004; // x = -19.9844, f(x) = 0.0000
    12'hB02: soft_out = 32'h00000005; // x = -19.9688, f(x) = 0.0000
    12'hB03: soft_out = 32'h00000005; // x = -19.9531, f(x) = 0.0000
    12'hB04: soft_out = 32'h00000005; // x = -19.9375, f(x) = 0.0000
    12'hB05: soft_out = 32'h00000005; // x = -19.9219, f(x) = 0.0000
    12'hB06: soft_out = 32'h00000005; // x = -19.9062, f(x) = 0.0000
    12'hB07: soft_out = 32'h00000005; // x = -19.8906, f(x) = 0.0000
    12'hB08: soft_out = 32'h00000005; // x = -19.8750, f(x) = 0.0000
    12'hB09: soft_out = 32'h00000005; // x = -19.8594, f(x) = 0.0000
    12'hB0A: soft_out = 32'h00000005; // x = -19.8438, f(x) = 0.0000
    12'hB0B: soft_out = 32'h00000005; // x = -19.8281, f(x) = 0.0000
    12'hB0C: soft_out = 32'h00000005; // x = -19.8125, f(x) = 0.0000
    12'hB0D: soft_out = 32'h00000005; // x = -19.7969, f(x) = 0.0000
    12'hB0E: soft_out = 32'h00000006; // x = -19.7812, f(x) = 0.0000
    12'hB0F: soft_out = 32'h00000006; // x = -19.7656, f(x) = 0.0000
    12'hB10: soft_out = 32'h00000006; // x = -19.7500, f(x) = 0.0000
    12'hB11: soft_out = 32'h00000006; // x = -19.7344, f(x) = 0.0000
    12'hB12: soft_out = 32'h00000006; // x = -19.7188, f(x) = 0.0000
    12'hB13: soft_out = 32'h00000006; // x = -19.7031, f(x) = 0.0000
    12'hB14: soft_out = 32'h00000006; // x = -19.6875, f(x) = 0.0000
    12'hB15: soft_out = 32'h00000006; // x = -19.6719, f(x) = 0.0000
    12'hB16: soft_out = 32'h00000006; // x = -19.6562, f(x) = 0.0000
    12'hB17: soft_out = 32'h00000006; // x = -19.6406, f(x) = 0.0000
    12'hB18: soft_out = 32'h00000006; // x = -19.6250, f(x) = 0.0000
    12'hB19: soft_out = 32'h00000007; // x = -19.6094, f(x) = 0.0000
    12'hB1A: soft_out = 32'h00000007; // x = -19.5938, f(x) = 0.0000
    12'hB1B: soft_out = 32'h00000007; // x = -19.5781, f(x) = 0.0000
    12'hB1C: soft_out = 32'h00000007; // x = -19.5625, f(x) = 0.0000
    12'hB1D: soft_out = 32'h00000007; // x = -19.5469, f(x) = 0.0000
    12'hB1E: soft_out = 32'h00000007; // x = -19.5312, f(x) = 0.0000
    12'hB1F: soft_out = 32'h00000007; // x = -19.5156, f(x) = 0.0000
    12'hB20: soft_out = 32'h00000007; // x = -19.5000, f(x) = 0.0000
    12'hB21: soft_out = 32'h00000007; // x = -19.4844, f(x) = 0.0000
    12'hB22: soft_out = 32'h00000008; // x = -19.4688, f(x) = 0.0000
    12'hB23: soft_out = 32'h00000008; // x = -19.4531, f(x) = 0.0000
    12'hB24: soft_out = 32'h00000008; // x = -19.4375, f(x) = 0.0000
    12'hB25: soft_out = 32'h00000008; // x = -19.4219, f(x) = 0.0000
    12'hB26: soft_out = 32'h00000008; // x = -19.4062, f(x) = 0.0000
    12'hB27: soft_out = 32'h00000008; // x = -19.3906, f(x) = 0.0000
    12'hB28: soft_out = 32'h00000008; // x = -19.3750, f(x) = 0.0000
    12'hB29: soft_out = 32'h00000008; // x = -19.3594, f(x) = 0.0000
    12'hB2A: soft_out = 32'h00000009; // x = -19.3438, f(x) = 0.0000
    12'hB2B: soft_out = 32'h00000009; // x = -19.3281, f(x) = 0.0000
    12'hB2C: soft_out = 32'h00000009; // x = -19.3125, f(x) = 0.0000
    12'hB2D: soft_out = 32'h00000009; // x = -19.2969, f(x) = 0.0000
    12'hB2E: soft_out = 32'h00000009; // x = -19.2812, f(x) = 0.0000
    12'hB2F: soft_out = 32'h00000009; // x = -19.2656, f(x) = 0.0000
    12'hB30: soft_out = 32'h00000009; // x = -19.2500, f(x) = 0.0000
    12'hB31: soft_out = 32'h0000000A; // x = -19.2344, f(x) = 0.0000
    12'hB32: soft_out = 32'h0000000A; // x = -19.2188, f(x) = 0.0000
    12'hB33: soft_out = 32'h0000000A; // x = -19.2031, f(x) = 0.0000
    12'hB34: soft_out = 32'h0000000A; // x = -19.1875, f(x) = 0.0000
    12'hB35: soft_out = 32'h0000000A; // x = -19.1719, f(x) = 0.0000
    12'hB36: soft_out = 32'h0000000A; // x = -19.1562, f(x) = 0.0000
    12'hB37: soft_out = 32'h0000000A; // x = -19.1406, f(x) = 0.0000
    12'hB38: soft_out = 32'h0000000B; // x = -19.1250, f(x) = 0.0000
    12'hB39: soft_out = 32'h0000000B; // x = -19.1094, f(x) = 0.0000
    12'hB3A: soft_out = 32'h0000000B; // x = -19.0938, f(x) = 0.0000
    12'hB3B: soft_out = 32'h0000000B; // x = -19.0781, f(x) = 0.0000
    12'hB3C: soft_out = 32'h0000000B; // x = -19.0625, f(x) = 0.0000
    12'hB3D: soft_out = 32'h0000000B; // x = -19.0469, f(x) = 0.0000
    12'hB3E: soft_out = 32'h0000000C; // x = -19.0312, f(x) = 0.0000
    12'hB3F: soft_out = 32'h0000000C; // x = -19.0156, f(x) = 0.0000
    12'hB40: soft_out = 32'h0000000C; // x = -19.0000, f(x) = 0.0000
    12'hB41: soft_out = 32'h0000000C; // x = -18.9844, f(x) = 0.0000
    12'hB42: soft_out = 32'h0000000C; // x = -18.9688, f(x) = 0.0000
    12'hB43: soft_out = 32'h0000000D; // x = -18.9531, f(x) = 0.0000
    12'hB44: soft_out = 32'h0000000D; // x = -18.9375, f(x) = 0.0000
    12'hB45: soft_out = 32'h0000000D; // x = -18.9219, f(x) = 0.0000
    12'hB46: soft_out = 32'h0000000D; // x = -18.9062, f(x) = 0.0000
    12'hB47: soft_out = 32'h0000000D; // x = -18.8906, f(x) = 0.0000
    12'hB48: soft_out = 32'h0000000E; // x = -18.8750, f(x) = 0.0000
    12'hB49: soft_out = 32'h0000000E; // x = -18.8594, f(x) = 0.0000
    12'hB4A: soft_out = 32'h0000000E; // x = -18.8438, f(x) = 0.0000
    12'hB4B: soft_out = 32'h0000000E; // x = -18.8281, f(x) = 0.0000
    12'hB4C: soft_out = 32'h0000000F; // x = -18.8125, f(x) = 0.0000
    12'hB4D: soft_out = 32'h0000000F; // x = -18.7969, f(x) = 0.0000
    12'hB4E: soft_out = 32'h0000000F; // x = -18.7812, f(x) = 0.0000
    12'hB4F: soft_out = 32'h0000000F; // x = -18.7656, f(x) = 0.0000
    12'hB50: soft_out = 32'h0000000F; // x = -18.7500, f(x) = 0.0000
    12'hB51: soft_out = 32'h00000010; // x = -18.7344, f(x) = 0.0000
    12'hB52: soft_out = 32'h00000010; // x = -18.7188, f(x) = 0.0000
    12'hB53: soft_out = 32'h00000010; // x = -18.7031, f(x) = 0.0000
    12'hB54: soft_out = 32'h00000010; // x = -18.6875, f(x) = 0.0000
    12'hB55: soft_out = 32'h00000011; // x = -18.6719, f(x) = 0.0000
    12'hB56: soft_out = 32'h00000011; // x = -18.6562, f(x) = 0.0000
    12'hB57: soft_out = 32'h00000011; // x = -18.6406, f(x) = 0.0000
    12'hB58: soft_out = 32'h00000012; // x = -18.6250, f(x) = 0.0000
    12'hB59: soft_out = 32'h00000012; // x = -18.6094, f(x) = 0.0000
    12'hB5A: soft_out = 32'h00000012; // x = -18.5938, f(x) = 0.0000
    12'hB5B: soft_out = 32'h00000012; // x = -18.5781, f(x) = 0.0000
    12'hB5C: soft_out = 32'h00000013; // x = -18.5625, f(x) = 0.0000
    12'hB5D: soft_out = 32'h00000013; // x = -18.5469, f(x) = 0.0000
    12'hB5E: soft_out = 32'h00000013; // x = -18.5312, f(x) = 0.0000
    12'hB5F: soft_out = 32'h00000014; // x = -18.5156, f(x) = 0.0000
    12'hB60: soft_out = 32'h00000014; // x = -18.5000, f(x) = 0.0000
    12'hB61: soft_out = 32'h00000014; // x = -18.4844, f(x) = 0.0000
    12'hB62: soft_out = 32'h00000014; // x = -18.4688, f(x) = 0.0000
    12'hB63: soft_out = 32'h00000015; // x = -18.4531, f(x) = 0.0000
    12'hB64: soft_out = 32'h00000015; // x = -18.4375, f(x) = 0.0000
    12'hB65: soft_out = 32'h00000015; // x = -18.4219, f(x) = 0.0000
    12'hB66: soft_out = 32'h00000016; // x = -18.4062, f(x) = 0.0000
    12'hB67: soft_out = 32'h00000016; // x = -18.3906, f(x) = 0.0000
    12'hB68: soft_out = 32'h00000016; // x = -18.3750, f(x) = 0.0000
    12'hB69: soft_out = 32'h00000017; // x = -18.3594, f(x) = 0.0000
    12'hB6A: soft_out = 32'h00000017; // x = -18.3438, f(x) = 0.0000
    12'hB6B: soft_out = 32'h00000018; // x = -18.3281, f(x) = 0.0000
    12'hB6C: soft_out = 32'h00000018; // x = -18.3125, f(x) = 0.0000
    12'hB6D: soft_out = 32'h00000018; // x = -18.2969, f(x) = 0.0000
    12'hB6E: soft_out = 32'h00000019; // x = -18.2812, f(x) = 0.0000
    12'hB6F: soft_out = 32'h00000019; // x = -18.2656, f(x) = 0.0000
    12'hB70: soft_out = 32'h00000019; // x = -18.2500, f(x) = 0.0000
    12'hB71: soft_out = 32'h0000001A; // x = -18.2344, f(x) = 0.0000
    12'hB72: soft_out = 32'h0000001A; // x = -18.2188, f(x) = 0.0000
    12'hB73: soft_out = 32'h0000001B; // x = -18.2031, f(x) = 0.0000
    12'hB74: soft_out = 32'h0000001B; // x = -18.1875, f(x) = 0.0000
    12'hB75: soft_out = 32'h0000001C; // x = -18.1719, f(x) = 0.0000
    12'hB76: soft_out = 32'h0000001C; // x = -18.1562, f(x) = 0.0000
    12'hB77: soft_out = 32'h0000001C; // x = -18.1406, f(x) = 0.0000
    12'hB78: soft_out = 32'h0000001D; // x = -18.1250, f(x) = 0.0000
    12'hB79: soft_out = 32'h0000001D; // x = -18.1094, f(x) = 0.0000
    12'hB7A: soft_out = 32'h0000001E; // x = -18.0938, f(x) = 0.0000
    12'hB7B: soft_out = 32'h0000001E; // x = -18.0781, f(x) = 0.0000
    12'hB7C: soft_out = 32'h0000001F; // x = -18.0625, f(x) = 0.0000
    12'hB7D: soft_out = 32'h0000001F; // x = -18.0469, f(x) = 0.0000
    12'hB7E: soft_out = 32'h00000020; // x = -18.0312, f(x) = 0.0000
    12'hB7F: soft_out = 32'h00000020; // x = -18.0156, f(x) = 0.0000
    12'hB80: soft_out = 32'h00000021; // x = -18.0000, f(x) = 0.0000
    12'hB81: soft_out = 32'h00000021; // x = -17.9844, f(x) = 0.0000
    12'hB82: soft_out = 32'h00000022; // x = -17.9688, f(x) = 0.0000
    12'hB83: soft_out = 32'h00000022; // x = -17.9531, f(x) = 0.0000
    12'hB84: soft_out = 32'h00000023; // x = -17.9375, f(x) = 0.0000
    12'hB85: soft_out = 32'h00000023; // x = -17.9219, f(x) = 0.0000
    12'hB86: soft_out = 32'h00000024; // x = -17.9062, f(x) = 0.0000
    12'hB87: soft_out = 32'h00000024; // x = -17.8906, f(x) = 0.0000
    12'hB88: soft_out = 32'h00000025; // x = -17.8750, f(x) = 0.0000
    12'hB89: soft_out = 32'h00000026; // x = -17.8594, f(x) = 0.0000
    12'hB8A: soft_out = 32'h00000026; // x = -17.8438, f(x) = 0.0000
    12'hB8B: soft_out = 32'h00000027; // x = -17.8281, f(x) = 0.0000
    12'hB8C: soft_out = 32'h00000027; // x = -17.8125, f(x) = 0.0000
    12'hB8D: soft_out = 32'h00000028; // x = -17.7969, f(x) = 0.0000
    12'hB8E: soft_out = 32'h00000029; // x = -17.7812, f(x) = 0.0000
    12'hB8F: soft_out = 32'h00000029; // x = -17.7656, f(x) = 0.0000
    12'hB90: soft_out = 32'h0000002A; // x = -17.7500, f(x) = 0.0000
    12'hB91: soft_out = 32'h0000002B; // x = -17.7344, f(x) = 0.0000
    12'hB92: soft_out = 32'h0000002B; // x = -17.7188, f(x) = 0.0000
    12'hB93: soft_out = 32'h0000002C; // x = -17.7031, f(x) = 0.0000
    12'hB94: soft_out = 32'h0000002D; // x = -17.6875, f(x) = 0.0000
    12'hB95: soft_out = 32'h0000002D; // x = -17.6719, f(x) = 0.0000
    12'hB96: soft_out = 32'h0000002E; // x = -17.6562, f(x) = 0.0000
    12'hB97: soft_out = 32'h0000002F; // x = -17.6406, f(x) = 0.0000
    12'hB98: soft_out = 32'h00000030; // x = -17.6250, f(x) = 0.0000
    12'hB99: soft_out = 32'h00000030; // x = -17.6094, f(x) = 0.0000
    12'hB9A: soft_out = 32'h00000031; // x = -17.5938, f(x) = 0.0000
    12'hB9B: soft_out = 32'h00000032; // x = -17.5781, f(x) = 0.0000
    12'hB9C: soft_out = 32'h00000033; // x = -17.5625, f(x) = 0.0000
    12'hB9D: soft_out = 32'h00000033; // x = -17.5469, f(x) = 0.0000
    12'hB9E: soft_out = 32'h00000034; // x = -17.5312, f(x) = 0.0000
    12'hB9F: soft_out = 32'h00000035; // x = -17.5156, f(x) = 0.0000
    12'hBA0: soft_out = 32'h00000036; // x = -17.5000, f(x) = 0.0000
    12'hBA1: soft_out = 32'h00000037; // x = -17.4844, f(x) = 0.0000
    12'hBA2: soft_out = 32'h00000038; // x = -17.4688, f(x) = 0.0000
    12'hBA3: soft_out = 32'h00000039; // x = -17.4531, f(x) = 0.0000
    12'hBA4: soft_out = 32'h00000039; // x = -17.4375, f(x) = 0.0000
    12'hBA5: soft_out = 32'h0000003A; // x = -17.4219, f(x) = 0.0000
    12'hBA6: soft_out = 32'h0000003B; // x = -17.4062, f(x) = 0.0000
    12'hBA7: soft_out = 32'h0000003C; // x = -17.3906, f(x) = 0.0000
    12'hBA8: soft_out = 32'h0000003D; // x = -17.3750, f(x) = 0.0000
    12'hBA9: soft_out = 32'h0000003E; // x = -17.3594, f(x) = 0.0000
    12'hBAA: soft_out = 32'h0000003F; // x = -17.3438, f(x) = 0.0000
    12'hBAB: soft_out = 32'h00000040; // x = -17.3281, f(x) = 0.0000
    12'hBAC: soft_out = 32'h00000041; // x = -17.3125, f(x) = 0.0000
    12'hBAD: soft_out = 32'h00000042; // x = -17.2969, f(x) = 0.0000
    12'hBAE: soft_out = 32'h00000043; // x = -17.2812, f(x) = 0.0000
    12'hBAF: soft_out = 32'h00000044; // x = -17.2656, f(x) = 0.0000
    12'hBB0: soft_out = 32'h00000045; // x = -17.2500, f(x) = 0.0000
    12'hBB1: soft_out = 32'h00000046; // x = -17.2344, f(x) = 0.0000
    12'hBB2: soft_out = 32'h00000047; // x = -17.2188, f(x) = 0.0000
    12'hBB3: soft_out = 32'h00000049; // x = -17.2031, f(x) = 0.0000
    12'hBB4: soft_out = 32'h0000004A; // x = -17.1875, f(x) = 0.0000
    12'hBB5: soft_out = 32'h0000004B; // x = -17.1719, f(x) = 0.0000
    12'hBB6: soft_out = 32'h0000004C; // x = -17.1562, f(x) = 0.0000
    12'hBB7: soft_out = 32'h0000004D; // x = -17.1406, f(x) = 0.0000
    12'hBB8: soft_out = 32'h0000004E; // x = -17.1250, f(x) = 0.0000
    12'hBB9: soft_out = 32'h00000050; // x = -17.1094, f(x) = 0.0000
    12'hBBA: soft_out = 32'h00000051; // x = -17.0938, f(x) = 0.0000
    12'hBBB: soft_out = 32'h00000052; // x = -17.0781, f(x) = 0.0000
    12'hBBC: soft_out = 32'h00000054; // x = -17.0625, f(x) = 0.0000
    12'hBBD: soft_out = 32'h00000055; // x = -17.0469, f(x) = 0.0000
    12'hBBE: soft_out = 32'h00000056; // x = -17.0312, f(x) = 0.0000
    12'hBBF: soft_out = 32'h00000058; // x = -17.0156, f(x) = 0.0000
    12'hBC0: soft_out = 32'h00000059; // x = -17.0000, f(x) = 0.0000
    12'hBC1: soft_out = 32'h0000005A; // x = -16.9844, f(x) = 0.0000
    12'hBC2: soft_out = 32'h0000005C; // x = -16.9688, f(x) = 0.0000
    12'hBC3: soft_out = 32'h0000005D; // x = -16.9531, f(x) = 0.0000
    12'hBC4: soft_out = 32'h0000005F; // x = -16.9375, f(x) = 0.0000
    12'hBC5: soft_out = 32'h00000060; // x = -16.9219, f(x) = 0.0000
    12'hBC6: soft_out = 32'h00000062; // x = -16.9062, f(x) = 0.0000
    12'hBC7: soft_out = 32'h00000063; // x = -16.8906, f(x) = 0.0000
    12'hBC8: soft_out = 32'h00000065; // x = -16.8750, f(x) = 0.0000
    12'hBC9: soft_out = 32'h00000066; // x = -16.8594, f(x) = 0.0000
    12'hBCA: soft_out = 32'h00000068; // x = -16.8438, f(x) = 0.0000
    12'hBCB: soft_out = 32'h0000006A; // x = -16.8281, f(x) = 0.0000
    12'hBCC: soft_out = 32'h0000006B; // x = -16.8125, f(x) = 0.0000
    12'hBCD: soft_out = 32'h0000006D; // x = -16.7969, f(x) = 0.0000
    12'hBCE: soft_out = 32'h0000006F; // x = -16.7812, f(x) = 0.0000
    12'hBCF: soft_out = 32'h00000070; // x = -16.7656, f(x) = 0.0000
    12'hBD0: soft_out = 32'h00000072; // x = -16.7500, f(x) = 0.0000
    12'hBD1: soft_out = 32'h00000074; // x = -16.7344, f(x) = 0.0000
    12'hBD2: soft_out = 32'h00000076; // x = -16.7188, f(x) = 0.0000
    12'hBD3: soft_out = 32'h00000078; // x = -16.7031, f(x) = 0.0000
    12'hBD4: soft_out = 32'h0000007A; // x = -16.6875, f(x) = 0.0000
    12'hBD5: soft_out = 32'h0000007B; // x = -16.6719, f(x) = 0.0000
    12'hBD6: soft_out = 32'h0000007D; // x = -16.6562, f(x) = 0.0000
    12'hBD7: soft_out = 32'h0000007F; // x = -16.6406, f(x) = 0.0000
    12'hBD8: soft_out = 32'h00000081; // x = -16.6250, f(x) = 0.0000
    12'hBD9: soft_out = 32'h00000083; // x = -16.6094, f(x) = 0.0000
    12'hBDA: soft_out = 32'h00000085; // x = -16.5938, f(x) = 0.0000
    12'hBDB: soft_out = 32'h00000088; // x = -16.5781, f(x) = 0.0000
    12'hBDC: soft_out = 32'h0000008A; // x = -16.5625, f(x) = 0.0000
    12'hBDD: soft_out = 32'h0000008C; // x = -16.5469, f(x) = 0.0000
    12'hBDE: soft_out = 32'h0000008E; // x = -16.5312, f(x) = 0.0000
    12'hBDF: soft_out = 32'h00000090; // x = -16.5156, f(x) = 0.0000
    12'hBE0: soft_out = 32'h00000093; // x = -16.5000, f(x) = 0.0000
    12'hBE1: soft_out = 32'h00000095; // x = -16.4844, f(x) = 0.0000
    12'hBE2: soft_out = 32'h00000097; // x = -16.4688, f(x) = 0.0000
    12'hBE3: soft_out = 32'h0000009A; // x = -16.4531, f(x) = 0.0000
    12'hBE4: soft_out = 32'h0000009C; // x = -16.4375, f(x) = 0.0000
    12'hBE5: soft_out = 32'h0000009E; // x = -16.4219, f(x) = 0.0000
    12'hBE6: soft_out = 32'h000000A1; // x = -16.4062, f(x) = 0.0000
    12'hBE7: soft_out = 32'h000000A4; // x = -16.3906, f(x) = 0.0000
    12'hBE8: soft_out = 32'h000000A6; // x = -16.3750, f(x) = 0.0000
    12'hBE9: soft_out = 32'h000000A9; // x = -16.3594, f(x) = 0.0000
    12'hBEA: soft_out = 32'h000000AB; // x = -16.3438, f(x) = 0.0000
    12'hBEB: soft_out = 32'h000000AE; // x = -16.3281, f(x) = 0.0000
    12'hBEC: soft_out = 32'h000000B1; // x = -16.3125, f(x) = 0.0000
    12'hBED: soft_out = 32'h000000B4; // x = -16.2969, f(x) = 0.0000
    12'hBEE: soft_out = 32'h000000B6; // x = -16.2812, f(x) = 0.0000
    12'hBEF: soft_out = 32'h000000B9; // x = -16.2656, f(x) = 0.0000
    12'hBF0: soft_out = 32'h000000BC; // x = -16.2500, f(x) = 0.0000
    12'hBF1: soft_out = 32'h000000BF; // x = -16.2344, f(x) = 0.0000
    12'hBF2: soft_out = 32'h000000C2; // x = -16.2188, f(x) = 0.0000
    12'hBF3: soft_out = 32'h000000C5; // x = -16.2031, f(x) = 0.0000
    12'hBF4: soft_out = 32'h000000C8; // x = -16.1875, f(x) = 0.0000
    12'hBF5: soft_out = 32'h000000CC; // x = -16.1719, f(x) = 0.0000
    12'hBF6: soft_out = 32'h000000CF; // x = -16.1562, f(x) = 0.0000
    12'hBF7: soft_out = 32'h000000D2; // x = -16.1406, f(x) = 0.0000
    12'hBF8: soft_out = 32'h000000D5; // x = -16.1250, f(x) = 0.0000
    12'hBF9: soft_out = 32'h000000D9; // x = -16.1094, f(x) = 0.0000
    12'hBFA: soft_out = 32'h000000DC; // x = -16.0938, f(x) = 0.0000
    12'hBFB: soft_out = 32'h000000E0; // x = -16.0781, f(x) = 0.0000
    12'hBFC: soft_out = 32'h000000E3; // x = -16.0625, f(x) = 0.0000
    12'hBFD: soft_out = 32'h000000E7; // x = -16.0469, f(x) = 0.0000
    12'hBFE: soft_out = 32'h000000EA; // x = -16.0312, f(x) = 0.0000
    12'hBFF: soft_out = 32'h000000EE; // x = -16.0156, f(x) = 0.0000
    12'hC00: soft_out = 32'h000000F2; // x = -16.0000, f(x) = 0.0000
    12'hC01: soft_out = 32'h000000F5; // x = -15.9844, f(x) = 0.0000
    12'hC02: soft_out = 32'h000000F9; // x = -15.9688, f(x) = 0.0000
    12'hC03: soft_out = 32'h000000FD; // x = -15.9531, f(x) = 0.0000
    12'hC04: soft_out = 32'h00000101; // x = -15.9375, f(x) = 0.0000
    12'hC05: soft_out = 32'h00000105; // x = -15.9219, f(x) = 0.0000
    12'hC06: soft_out = 32'h00000109; // x = -15.9062, f(x) = 0.0000
    12'hC07: soft_out = 32'h0000010E; // x = -15.8906, f(x) = 0.0000
    12'hC08: soft_out = 32'h00000112; // x = -15.8750, f(x) = 0.0000
    12'hC09: soft_out = 32'h00000116; // x = -15.8594, f(x) = 0.0000
    12'hC0A: soft_out = 32'h0000011B; // x = -15.8438, f(x) = 0.0000
    12'hC0B: soft_out = 32'h0000011F; // x = -15.8281, f(x) = 0.0000
    12'hC0C: soft_out = 32'h00000124; // x = -15.8125, f(x) = 0.0000
    12'hC0D: soft_out = 32'h00000128; // x = -15.7969, f(x) = 0.0000
    12'hC0E: soft_out = 32'h0000012D; // x = -15.7812, f(x) = 0.0000
    12'hC0F: soft_out = 32'h00000131; // x = -15.7656, f(x) = 0.0000
    12'hC10: soft_out = 32'h00000136; // x = -15.7500, f(x) = 0.0000
    12'hC11: soft_out = 32'h0000013B; // x = -15.7344, f(x) = 0.0000
    12'hC12: soft_out = 32'h00000140; // x = -15.7188, f(x) = 0.0000
    12'hC13: soft_out = 32'h00000145; // x = -15.7031, f(x) = 0.0000
    12'hC14: soft_out = 32'h0000014A; // x = -15.6875, f(x) = 0.0000
    12'hC15: soft_out = 32'h00000150; // x = -15.6719, f(x) = 0.0000
    12'hC16: soft_out = 32'h00000155; // x = -15.6562, f(x) = 0.0000
    12'hC17: soft_out = 32'h0000015A; // x = -15.6406, f(x) = 0.0000
    12'hC18: soft_out = 32'h00000160; // x = -15.6250, f(x) = 0.0000
    12'hC19: soft_out = 32'h00000165; // x = -15.6094, f(x) = 0.0000
    12'hC1A: soft_out = 32'h0000016B; // x = -15.5938, f(x) = 0.0000
    12'hC1B: soft_out = 32'h00000170; // x = -15.5781, f(x) = 0.0000
    12'hC1C: soft_out = 32'h00000176; // x = -15.5625, f(x) = 0.0000
    12'hC1D: soft_out = 32'h0000017C; // x = -15.5469, f(x) = 0.0000
    12'hC1E: soft_out = 32'h00000182; // x = -15.5312, f(x) = 0.0000
    12'hC1F: soft_out = 32'h00000188; // x = -15.5156, f(x) = 0.0000
    12'hC20: soft_out = 32'h0000018E; // x = -15.5000, f(x) = 0.0000
    12'hC21: soft_out = 32'h00000195; // x = -15.4844, f(x) = 0.0000
    12'hC22: soft_out = 32'h0000019B; // x = -15.4688, f(x) = 0.0000
    12'hC23: soft_out = 32'h000001A2; // x = -15.4531, f(x) = 0.0000
    12'hC24: soft_out = 32'h000001A8; // x = -15.4375, f(x) = 0.0000
    12'hC25: soft_out = 32'h000001AF; // x = -15.4219, f(x) = 0.0000
    12'hC26: soft_out = 32'h000001B6; // x = -15.4062, f(x) = 0.0000
    12'hC27: soft_out = 32'h000001BC; // x = -15.3906, f(x) = 0.0000
    12'hC28: soft_out = 32'h000001C3; // x = -15.3750, f(x) = 0.0000
    12'hC29: soft_out = 32'h000001CB; // x = -15.3594, f(x) = 0.0000
    12'hC2A: soft_out = 32'h000001D2; // x = -15.3438, f(x) = 0.0000
    12'hC2B: soft_out = 32'h000001D9; // x = -15.3281, f(x) = 0.0000
    12'hC2C: soft_out = 32'h000001E1; // x = -15.3125, f(x) = 0.0000
    12'hC2D: soft_out = 32'h000001E8; // x = -15.2969, f(x) = 0.0000
    12'hC2E: soft_out = 32'h000001F0; // x = -15.2812, f(x) = 0.0000
    12'hC2F: soft_out = 32'h000001F8; // x = -15.2656, f(x) = 0.0000
    12'hC30: soft_out = 32'h00000200; // x = -15.2500, f(x) = 0.0000
    12'hC31: soft_out = 32'h00000208; // x = -15.2344, f(x) = 0.0000
    12'hC32: soft_out = 32'h00000210; // x = -15.2188, f(x) = 0.0000
    12'hC33: soft_out = 32'h00000218; // x = -15.2031, f(x) = 0.0000
    12'hC34: soft_out = 32'h00000221; // x = -15.1875, f(x) = 0.0000
    12'hC35: soft_out = 32'h00000229; // x = -15.1719, f(x) = 0.0000
    12'hC36: soft_out = 32'h00000232; // x = -15.1562, f(x) = 0.0000
    12'hC37: soft_out = 32'h0000023B; // x = -15.1406, f(x) = 0.0000
    12'hC38: soft_out = 32'h00000244; // x = -15.1250, f(x) = 0.0000
    12'hC39: soft_out = 32'h0000024D; // x = -15.1094, f(x) = 0.0000
    12'hC3A: soft_out = 32'h00000256; // x = -15.0938, f(x) = 0.0000
    12'hC3B: soft_out = 32'h00000260; // x = -15.0781, f(x) = 0.0000
    12'hC3C: soft_out = 32'h00000269; // x = -15.0625, f(x) = 0.0000
    12'hC3D: soft_out = 32'h00000273; // x = -15.0469, f(x) = 0.0000
    12'hC3E: soft_out = 32'h0000027D; // x = -15.0312, f(x) = 0.0000
    12'hC3F: soft_out = 32'h00000287; // x = -15.0156, f(x) = 0.0000
    12'hC40: soft_out = 32'h00000291; // x = -15.0000, f(x) = 0.0000
    12'hC41: soft_out = 32'h0000029B; // x = -14.9844, f(x) = 0.0000
    12'hC42: soft_out = 32'h000002A6; // x = -14.9688, f(x) = 0.0000
    12'hC43: soft_out = 32'h000002B0; // x = -14.9531, f(x) = 0.0000
    12'hC44: soft_out = 32'h000002BB; // x = -14.9375, f(x) = 0.0000
    12'hC45: soft_out = 32'h000002C6; // x = -14.9219, f(x) = 0.0000
    12'hC46: soft_out = 32'h000002D1; // x = -14.9062, f(x) = 0.0000
    12'hC47: soft_out = 32'h000002DD; // x = -14.8906, f(x) = 0.0000
    12'hC48: soft_out = 32'h000002E8; // x = -14.8750, f(x) = 0.0000
    12'hC49: soft_out = 32'h000002F4; // x = -14.8594, f(x) = 0.0000
    12'hC4A: soft_out = 32'h00000300; // x = -14.8438, f(x) = 0.0000
    12'hC4B: soft_out = 32'h0000030C; // x = -14.8281, f(x) = 0.0000
    12'hC4C: soft_out = 32'h00000318; // x = -14.8125, f(x) = 0.0000
    12'hC4D: soft_out = 32'h00000325; // x = -14.7969, f(x) = 0.0000
    12'hC4E: soft_out = 32'h00000332; // x = -14.7812, f(x) = 0.0000
    12'hC4F: soft_out = 32'h0000033E; // x = -14.7656, f(x) = 0.0000
    12'hC50: soft_out = 32'h0000034C; // x = -14.7500, f(x) = 0.0000
    12'hC51: soft_out = 32'h00000359; // x = -14.7344, f(x) = 0.0000
    12'hC52: soft_out = 32'h00000366; // x = -14.7188, f(x) = 0.0000
    12'hC53: soft_out = 32'h00000374; // x = -14.7031, f(x) = 0.0000
    12'hC54: soft_out = 32'h00000382; // x = -14.6875, f(x) = 0.0000
    12'hC55: soft_out = 32'h00000390; // x = -14.6719, f(x) = 0.0000
    12'hC56: soft_out = 32'h0000039E; // x = -14.6562, f(x) = 0.0000
    12'hC57: soft_out = 32'h000003AD; // x = -14.6406, f(x) = 0.0000
    12'hC58: soft_out = 32'h000003BC; // x = -14.6250, f(x) = 0.0000
    12'hC59: soft_out = 32'h000003CB; // x = -14.6094, f(x) = 0.0000
    12'hC5A: soft_out = 32'h000003DA; // x = -14.5938, f(x) = 0.0000
    12'hC5B: soft_out = 32'h000003EA; // x = -14.5781, f(x) = 0.0000
    12'hC5C: soft_out = 32'h000003F9; // x = -14.5625, f(x) = 0.0000
    12'hC5D: soft_out = 32'h00000409; // x = -14.5469, f(x) = 0.0000
    12'hC5E: soft_out = 32'h0000041A; // x = -14.5312, f(x) = 0.0000
    12'hC5F: soft_out = 32'h0000042A; // x = -14.5156, f(x) = 0.0000
    12'hC60: soft_out = 32'h0000043B; // x = -14.5000, f(x) = 0.0000
    12'hC61: soft_out = 32'h0000044C; // x = -14.4844, f(x) = 0.0000
    12'hC62: soft_out = 32'h0000045D; // x = -14.4688, f(x) = 0.0000
    12'hC63: soft_out = 32'h0000046F; // x = -14.4531, f(x) = 0.0000
    12'hC64: soft_out = 32'h00000481; // x = -14.4375, f(x) = 0.0000
    12'hC65: soft_out = 32'h00000493; // x = -14.4219, f(x) = 0.0000
    12'hC66: soft_out = 32'h000004A6; // x = -14.4062, f(x) = 0.0000
    12'hC67: soft_out = 32'h000004B8; // x = -14.3906, f(x) = 0.0000
    12'hC68: soft_out = 32'h000004CB; // x = -14.3750, f(x) = 0.0000
    12'hC69: soft_out = 32'h000004DF; // x = -14.3594, f(x) = 0.0000
    12'hC6A: soft_out = 32'h000004F2; // x = -14.3438, f(x) = 0.0000
    12'hC6B: soft_out = 32'h00000506; // x = -14.3281, f(x) = 0.0000
    12'hC6C: soft_out = 32'h0000051A; // x = -14.3125, f(x) = 0.0000
    12'hC6D: soft_out = 32'h0000052F; // x = -14.2969, f(x) = 0.0000
    12'hC6E: soft_out = 32'h00000544; // x = -14.2812, f(x) = 0.0000
    12'hC6F: soft_out = 32'h00000559; // x = -14.2656, f(x) = 0.0000
    12'hC70: soft_out = 32'h0000056F; // x = -14.2500, f(x) = 0.0000
    12'hC71: soft_out = 32'h00000585; // x = -14.2344, f(x) = 0.0000
    12'hC72: soft_out = 32'h0000059B; // x = -14.2188, f(x) = 0.0000
    12'hC73: soft_out = 32'h000005B1; // x = -14.2031, f(x) = 0.0000
    12'hC74: soft_out = 32'h000005C8; // x = -14.1875, f(x) = 0.0000
    12'hC75: soft_out = 32'h000005E0; // x = -14.1719, f(x) = 0.0000
    12'hC76: soft_out = 32'h000005F7; // x = -14.1562, f(x) = 0.0000
    12'hC77: soft_out = 32'h0000060F; // x = -14.1406, f(x) = 0.0000
    12'hC78: soft_out = 32'h00000628; // x = -14.1250, f(x) = 0.0000
    12'hC79: soft_out = 32'h00000641; // x = -14.1094, f(x) = 0.0000
    12'hC7A: soft_out = 32'h0000065A; // x = -14.0938, f(x) = 0.0000
    12'hC7B: soft_out = 32'h00000673; // x = -14.0781, f(x) = 0.0000
    12'hC7C: soft_out = 32'h0000068E; // x = -14.0625, f(x) = 0.0000
    12'hC7D: soft_out = 32'h000006A8; // x = -14.0469, f(x) = 0.0000
    12'hC7E: soft_out = 32'h000006C3; // x = -14.0312, f(x) = 0.0000
    12'hC7F: soft_out = 32'h000006DE; // x = -14.0156, f(x) = 0.0000
    12'hC80: soft_out = 32'h000006FA; // x = -14.0000, f(x) = 0.0000
    12'hC81: soft_out = 32'h00000716; // x = -13.9844, f(x) = 0.0000
    12'hC82: soft_out = 32'h00000732; // x = -13.9688, f(x) = 0.0000
    12'hC83: soft_out = 32'h0000074F; // x = -13.9531, f(x) = 0.0000
    12'hC84: soft_out = 32'h0000076D; // x = -13.9375, f(x) = 0.0000
    12'hC85: soft_out = 32'h0000078B; // x = -13.9219, f(x) = 0.0000
    12'hC86: soft_out = 32'h000007A9; // x = -13.9062, f(x) = 0.0000
    12'hC87: soft_out = 32'h000007C8; // x = -13.8906, f(x) = 0.0000
    12'hC88: soft_out = 32'h000007E7; // x = -13.8750, f(x) = 0.0000
    12'hC89: soft_out = 32'h00000807; // x = -13.8594, f(x) = 0.0000
    12'hC8A: soft_out = 32'h00000828; // x = -13.8438, f(x) = 0.0000
    12'hC8B: soft_out = 32'h00000849; // x = -13.8281, f(x) = 0.0000
    12'hC8C: soft_out = 32'h0000086A; // x = -13.8125, f(x) = 0.0000
    12'hC8D: soft_out = 32'h0000088C; // x = -13.7969, f(x) = 0.0000
    12'hC8E: soft_out = 32'h000008AE; // x = -13.7812, f(x) = 0.0000
    12'hC8F: soft_out = 32'h000008D1; // x = -13.7656, f(x) = 0.0000
    12'hC90: soft_out = 32'h000008F5; // x = -13.7500, f(x) = 0.0000
    12'hC91: soft_out = 32'h00000919; // x = -13.7344, f(x) = 0.0000
    12'hC92: soft_out = 32'h0000093E; // x = -13.7188, f(x) = 0.0000
    12'hC93: soft_out = 32'h00000963; // x = -13.7031, f(x) = 0.0000
    12'hC94: soft_out = 32'h00000989; // x = -13.6875, f(x) = 0.0000
    12'hC95: soft_out = 32'h000009AF; // x = -13.6719, f(x) = 0.0000
    12'hC96: soft_out = 32'h000009D6; // x = -13.6562, f(x) = 0.0000
    12'hC97: soft_out = 32'h000009FE; // x = -13.6406, f(x) = 0.0000
    12'hC98: soft_out = 32'h00000A26; // x = -13.6250, f(x) = 0.0000
    12'hC99: soft_out = 32'h00000A4F; // x = -13.6094, f(x) = 0.0000
    12'hC9A: soft_out = 32'h00000A79; // x = -13.5938, f(x) = 0.0000
    12'hC9B: soft_out = 32'h00000AA3; // x = -13.5781, f(x) = 0.0000
    12'hC9C: soft_out = 32'h00000ACE; // x = -13.5625, f(x) = 0.0000
    12'hC9D: soft_out = 32'h00000AF9; // x = -13.5469, f(x) = 0.0000
    12'hC9E: soft_out = 32'h00000B26; // x = -13.5312, f(x) = 0.0000
    12'hC9F: soft_out = 32'h00000B52; // x = -13.5156, f(x) = 0.0000
    12'hCA0: soft_out = 32'h00000B80; // x = -13.5000, f(x) = 0.0000
    12'hCA1: soft_out = 32'h00000BAE; // x = -13.4844, f(x) = 0.0000
    12'hCA2: soft_out = 32'h00000BDE; // x = -13.4688, f(x) = 0.0000
    12'hCA3: soft_out = 32'h00000C0D; // x = -13.4531, f(x) = 0.0000
    12'hCA4: soft_out = 32'h00000C3E; // x = -13.4375, f(x) = 0.0000
    12'hCA5: soft_out = 32'h00000C6F; // x = -13.4219, f(x) = 0.0000
    12'hCA6: soft_out = 32'h00000CA1; // x = -13.4062, f(x) = 0.0000
    12'hCA7: soft_out = 32'h00000CD4; // x = -13.3906, f(x) = 0.0000
    12'hCA8: soft_out = 32'h00000D08; // x = -13.3750, f(x) = 0.0000
    12'hCA9: soft_out = 32'h00000D3D; // x = -13.3594, f(x) = 0.0000
    12'hCAA: soft_out = 32'h00000D72; // x = -13.3438, f(x) = 0.0000
    12'hCAB: soft_out = 32'h00000DA8; // x = -13.3281, f(x) = 0.0000
    12'hCAC: soft_out = 32'h00000DDF; // x = -13.3125, f(x) = 0.0000
    12'hCAD: soft_out = 32'h00000E17; // x = -13.2969, f(x) = 0.0000
    12'hCAE: soft_out = 32'h00000E50; // x = -13.2812, f(x) = 0.0000
    12'hCAF: soft_out = 32'h00000E8A; // x = -13.2656, f(x) = 0.0000
    12'hCB0: soft_out = 32'h00000EC4; // x = -13.2500, f(x) = 0.0000
    12'hCB1: soft_out = 32'h00000F00; // x = -13.2344, f(x) = 0.0000
    12'hCB2: soft_out = 32'h00000F3C; // x = -13.2188, f(x) = 0.0000
    12'hCB3: soft_out = 32'h00000F7A; // x = -13.2031, f(x) = 0.0000
    12'hCB4: soft_out = 32'h00000FB8; // x = -13.1875, f(x) = 0.0000
    12'hCB5: soft_out = 32'h00000FF7; // x = -13.1719, f(x) = 0.0000
    12'hCB6: soft_out = 32'h00001038; // x = -13.1562, f(x) = 0.0000
    12'hCB7: soft_out = 32'h00001079; // x = -13.1406, f(x) = 0.0000
    12'hCB8: soft_out = 32'h000010BC; // x = -13.1250, f(x) = 0.0000
    12'hCB9: soft_out = 32'h000010FF; // x = -13.1094, f(x) = 0.0000
    12'hCBA: soft_out = 32'h00001144; // x = -13.0938, f(x) = 0.0000
    12'hCBB: soft_out = 32'h00001189; // x = -13.0781, f(x) = 0.0000
    12'hCBC: soft_out = 32'h000011D0; // x = -13.0625, f(x) = 0.0000
    12'hCBD: soft_out = 32'h00001218; // x = -13.0469, f(x) = 0.0000
    12'hCBE: soft_out = 32'h00001261; // x = -13.0312, f(x) = 0.0000
    12'hCBF: soft_out = 32'h000012AB; // x = -13.0156, f(x) = 0.0000
    12'hCC0: soft_out = 32'h000012F6; // x = -13.0000, f(x) = 0.0000
    12'hCC1: soft_out = 32'h00001342; // x = -12.9844, f(x) = 0.0000
    12'hCC2: soft_out = 32'h00001390; // x = -12.9688, f(x) = 0.0000
    12'hCC3: soft_out = 32'h000013DF; // x = -12.9531, f(x) = 0.0000
    12'hCC4: soft_out = 32'h0000142F; // x = -12.9375, f(x) = 0.0000
    12'hCC5: soft_out = 32'h00001480; // x = -12.9219, f(x) = 0.0000
    12'hCC6: soft_out = 32'h000014D3; // x = -12.9062, f(x) = 0.0000
    12'hCC7: soft_out = 32'h00001527; // x = -12.8906, f(x) = 0.0000
    12'hCC8: soft_out = 32'h0000157C; // x = -12.8750, f(x) = 0.0000
    12'hCC9: soft_out = 32'h000015D3; // x = -12.8594, f(x) = 0.0000
    12'hCCA: soft_out = 32'h0000162B; // x = -12.8438, f(x) = 0.0000
    12'hCCB: soft_out = 32'h00001684; // x = -12.8281, f(x) = 0.0000
    12'hCCC: soft_out = 32'h000016DF; // x = -12.8125, f(x) = 0.0000
    12'hCCD: soft_out = 32'h0000173B; // x = -12.7969, f(x) = 0.0000
    12'hCCE: soft_out = 32'h00001799; // x = -12.7812, f(x) = 0.0000
    12'hCCF: soft_out = 32'h000017F8; // x = -12.7656, f(x) = 0.0000
    12'hCD0: soft_out = 32'h00001859; // x = -12.7500, f(x) = 0.0000
    12'hCD1: soft_out = 32'h000018BB; // x = -12.7344, f(x) = 0.0000
    12'hCD2: soft_out = 32'h0000191F; // x = -12.7188, f(x) = 0.0000
    12'hCD3: soft_out = 32'h00001984; // x = -12.7031, f(x) = 0.0000
    12'hCD4: soft_out = 32'h000019EB; // x = -12.6875, f(x) = 0.0000
    12'hCD5: soft_out = 32'h00001A53; // x = -12.6719, f(x) = 0.0000
    12'hCD6: soft_out = 32'h00001ABD; // x = -12.6562, f(x) = 0.0000
    12'hCD7: soft_out = 32'h00001B29; // x = -12.6406, f(x) = 0.0000
    12'hCD8: soft_out = 32'h00001B97; // x = -12.6250, f(x) = 0.0000
    12'hCD9: soft_out = 32'h00001C06; // x = -12.6094, f(x) = 0.0000
    12'hCDA: soft_out = 32'h00001C77; // x = -12.5938, f(x) = 0.0000
    12'hCDB: soft_out = 32'h00001CE9; // x = -12.5781, f(x) = 0.0000
    12'hCDC: soft_out = 32'h00001D5E; // x = -12.5625, f(x) = 0.0000
    12'hCDD: soft_out = 32'h00001DD4; // x = -12.5469, f(x) = 0.0000
    12'hCDE: soft_out = 32'h00001E4D; // x = -12.5312, f(x) = 0.0000
    12'hCDF: soft_out = 32'h00001EC7; // x = -12.5156, f(x) = 0.0000
    12'hCE0: soft_out = 32'h00001F43; // x = -12.5000, f(x) = 0.0000
    12'hCE1: soft_out = 32'h00001FC1; // x = -12.4844, f(x) = 0.0000
    12'hCE2: soft_out = 32'h00002041; // x = -12.4688, f(x) = 0.0000
    12'hCE3: soft_out = 32'h000020C3; // x = -12.4531, f(x) = 0.0000
    12'hCE4: soft_out = 32'h00002147; // x = -12.4375, f(x) = 0.0000
    12'hCE5: soft_out = 32'h000021CD; // x = -12.4219, f(x) = 0.0000
    12'hCE6: soft_out = 32'h00002255; // x = -12.4062, f(x) = 0.0000
    12'hCE7: soft_out = 32'h000022E0; // x = -12.3906, f(x) = 0.0000
    12'hCE8: soft_out = 32'h0000236D; // x = -12.3750, f(x) = 0.0000
    12'hCE9: soft_out = 32'h000023FB; // x = -12.3594, f(x) = 0.0000
    12'hCEA: soft_out = 32'h0000248C; // x = -12.3438, f(x) = 0.0000
    12'hCEB: soft_out = 32'h00002520; // x = -12.3281, f(x) = 0.0000
    12'hCEC: soft_out = 32'h000025B5; // x = -12.3125, f(x) = 0.0000
    12'hCED: soft_out = 32'h0000264D; // x = -12.2969, f(x) = 0.0000
    12'hCEE: soft_out = 32'h000026E8; // x = -12.2812, f(x) = 0.0000
    12'hCEF: soft_out = 32'h00002785; // x = -12.2656, f(x) = 0.0000
    12'hCF0: soft_out = 32'h00002824; // x = -12.2500, f(x) = 0.0000
    12'hCF1: soft_out = 32'h000028C6; // x = -12.2344, f(x) = 0.0000
    12'hCF2: soft_out = 32'h0000296A; // x = -12.2188, f(x) = 0.0000
    12'hCF3: soft_out = 32'h00002A11; // x = -12.2031, f(x) = 0.0000
    12'hCF4: soft_out = 32'h00002ABB; // x = -12.1875, f(x) = 0.0000
    12'hCF5: soft_out = 32'h00002B67; // x = -12.1719, f(x) = 0.0000
    12'hCF6: soft_out = 32'h00002C16; // x = -12.1562, f(x) = 0.0000
    12'hCF7: soft_out = 32'h00002CC8; // x = -12.1406, f(x) = 0.0000
    12'hCF8: soft_out = 32'h00002D7C; // x = -12.1250, f(x) = 0.0000
    12'hCF9: soft_out = 32'h00002E34; // x = -12.1094, f(x) = 0.0000
    12'hCFA: soft_out = 32'h00002EEE; // x = -12.0938, f(x) = 0.0000
    12'hCFB: soft_out = 32'h00002FAB; // x = -12.0781, f(x) = 0.0000
    12'hCFC: soft_out = 32'h0000306B; // x = -12.0625, f(x) = 0.0000
    12'hCFD: soft_out = 32'h0000312E; // x = -12.0469, f(x) = 0.0000
    12'hCFE: soft_out = 32'h000031F5; // x = -12.0312, f(x) = 0.0000
    12'hCFF: soft_out = 32'h000032BE; // x = -12.0156, f(x) = 0.0000
    12'hD00: soft_out = 32'h0000338B; // x = -12.0000, f(x) = 0.0000
    12'hD01: soft_out = 32'h0000345A; // x = -11.9844, f(x) = 0.0000
    12'hD02: soft_out = 32'h0000352D; // x = -11.9688, f(x) = 0.0000
    12'hD03: soft_out = 32'h00003604; // x = -11.9531, f(x) = 0.0000
    12'hD04: soft_out = 32'h000036DE; // x = -11.9375, f(x) = 0.0000
    12'hD05: soft_out = 32'h000037BB; // x = -11.9219, f(x) = 0.0000
    12'hD06: soft_out = 32'h0000389B; // x = -11.9062, f(x) = 0.0000
    12'hD07: soft_out = 32'h00003980; // x = -11.8906, f(x) = 0.0000
    12'hD08: soft_out = 32'h00003A67; // x = -11.8750, f(x) = 0.0000
    12'hD09: soft_out = 32'h00003B53; // x = -11.8594, f(x) = 0.0000
    12'hD0A: soft_out = 32'h00003C42; // x = -11.8438, f(x) = 0.0000
    12'hD0B: soft_out = 32'h00003D35; // x = -11.8281, f(x) = 0.0000
    12'hD0C: soft_out = 32'h00003E2C; // x = -11.8125, f(x) = 0.0000
    12'hD0D: soft_out = 32'h00003F26; // x = -11.7969, f(x) = 0.0000
    12'hD0E: soft_out = 32'h00004025; // x = -11.7812, f(x) = 0.0000
    12'hD0F: soft_out = 32'h00004128; // x = -11.7656, f(x) = 0.0000
    12'hD10: soft_out = 32'h0000422E; // x = -11.7500, f(x) = 0.0000
    12'hD11: soft_out = 32'h00004339; // x = -11.7344, f(x) = 0.0000
    12'hD12: soft_out = 32'h00004448; // x = -11.7188, f(x) = 0.0000
    12'hD13: soft_out = 32'h0000455B; // x = -11.7031, f(x) = 0.0000
    12'hD14: soft_out = 32'h00004673; // x = -11.6875, f(x) = 0.0000
    12'hD15: soft_out = 32'h0000478F; // x = -11.6719, f(x) = 0.0000
    12'hD16: soft_out = 32'h000048AF; // x = -11.6562, f(x) = 0.0000
    12'hD17: soft_out = 32'h000049D4; // x = -11.6406, f(x) = 0.0000
    12'hD18: soft_out = 32'h00004AFE; // x = -11.6250, f(x) = 0.0000
    12'hD19: soft_out = 32'h00004C2C; // x = -11.6094, f(x) = 0.0000
    12'hD1A: soft_out = 32'h00004D5F; // x = -11.5938, f(x) = 0.0000
    12'hD1B: soft_out = 32'h00004E97; // x = -11.5781, f(x) = 0.0000
    12'hD1C: soft_out = 32'h00004FD4; // x = -11.5625, f(x) = 0.0000
    12'hD1D: soft_out = 32'h00005116; // x = -11.5469, f(x) = 0.0000
    12'hD1E: soft_out = 32'h0000525D; // x = -11.5312, f(x) = 0.0000
    12'hD1F: soft_out = 32'h000053A9; // x = -11.5156, f(x) = 0.0000
    12'hD20: soft_out = 32'h000054FA; // x = -11.5000, f(x) = 0.0000
    12'hD21: soft_out = 32'h00005651; // x = -11.4844, f(x) = 0.0000
    12'hD22: soft_out = 32'h000057AD; // x = -11.4688, f(x) = 0.0000
    12'hD23: soft_out = 32'h0000590E; // x = -11.4531, f(x) = 0.0000
    12'hD24: soft_out = 32'h00005A75; // x = -11.4375, f(x) = 0.0000
    12'hD25: soft_out = 32'h00005BE2; // x = -11.4219, f(x) = 0.0000
    12'hD26: soft_out = 32'h00005D54; // x = -11.4062, f(x) = 0.0000
    12'hD27: soft_out = 32'h00005ECD; // x = -11.3906, f(x) = 0.0000
    12'hD28: soft_out = 32'h0000604B; // x = -11.3750, f(x) = 0.0000
    12'hD29: soft_out = 32'h000061CF; // x = -11.3594, f(x) = 0.0000
    12'hD2A: soft_out = 32'h00006359; // x = -11.3438, f(x) = 0.0000
    12'hD2B: soft_out = 32'h000064EA; // x = -11.3281, f(x) = 0.0000
    12'hD2C: soft_out = 32'h00006681; // x = -11.3125, f(x) = 0.0000
    12'hD2D: soft_out = 32'h0000681E; // x = -11.2969, f(x) = 0.0000
    12'hD2E: soft_out = 32'h000069C2; // x = -11.2812, f(x) = 0.0000
    12'hD2F: soft_out = 32'h00006B6C; // x = -11.2656, f(x) = 0.0000
    12'hD30: soft_out = 32'h00006D1D; // x = -11.2500, f(x) = 0.0000
    12'hD31: soft_out = 32'h00006ED5; // x = -11.2344, f(x) = 0.0000
    12'hD32: soft_out = 32'h00007094; // x = -11.2188, f(x) = 0.0000
    12'hD33: soft_out = 32'h00007259; // x = -11.2031, f(x) = 0.0000
    12'hD34: soft_out = 32'h00007426; // x = -11.1875, f(x) = 0.0000
    12'hD35: soft_out = 32'h000075FB; // x = -11.1719, f(x) = 0.0000
    12'hD36: soft_out = 32'h000077D6; // x = -11.1562, f(x) = 0.0000
    12'hD37: soft_out = 32'h000079B9; // x = -11.1406, f(x) = 0.0000
    12'hD38: soft_out = 32'h00007BA4; // x = -11.1250, f(x) = 0.0000
    12'hD39: soft_out = 32'h00007D97; // x = -11.1094, f(x) = 0.0000
    12'hD3A: soft_out = 32'h00007F91; // x = -11.0938, f(x) = 0.0000
    12'hD3B: soft_out = 32'h00008193; // x = -11.0781, f(x) = 0.0000
    12'hD3C: soft_out = 32'h0000839E; // x = -11.0625, f(x) = 0.0000
    12'hD3D: soft_out = 32'h000085B0; // x = -11.0469, f(x) = 0.0000
    12'hD3E: soft_out = 32'h000087CB; // x = -11.0312, f(x) = 0.0000
    12'hD3F: soft_out = 32'h000089EF; // x = -11.0156, f(x) = 0.0000
    12'hD40: soft_out = 32'h00008C1B; // x = -11.0000, f(x) = 0.0000
    12'hD41: soft_out = 32'h00008E4F; // x = -10.9844, f(x) = 0.0000
    12'hD42: soft_out = 32'h0000908D; // x = -10.9688, f(x) = 0.0000
    12'hD43: soft_out = 32'h000092D4; // x = -10.9531, f(x) = 0.0000
    12'hD44: soft_out = 32'h00009524; // x = -10.9375, f(x) = 0.0000
    12'hD45: soft_out = 32'h0000977D; // x = -10.9219, f(x) = 0.0000
    12'hD46: soft_out = 32'h000099E0; // x = -10.9062, f(x) = 0.0000
    12'hD47: soft_out = 32'h00009C4C; // x = -10.8906, f(x) = 0.0000
    12'hD48: soft_out = 32'h00009EC2; // x = -10.8750, f(x) = 0.0000
    12'hD49: soft_out = 32'h0000A142; // x = -10.8594, f(x) = 0.0000
    12'hD4A: soft_out = 32'h0000A3CC; // x = -10.8438, f(x) = 0.0000
    12'hD4B: soft_out = 32'h0000A661; // x = -10.8281, f(x) = 0.0000
    12'hD4C: soft_out = 32'h0000A8FF; // x = -10.8125, f(x) = 0.0000
    12'hD4D: soft_out = 32'h0000ABA9; // x = -10.7969, f(x) = 0.0000
    12'hD4E: soft_out = 32'h0000AE5D; // x = -10.7812, f(x) = 0.0000
    12'hD4F: soft_out = 32'h0000B11C; // x = -10.7656, f(x) = 0.0000
    12'hD50: soft_out = 32'h0000B3E6; // x = -10.7500, f(x) = 0.0000
    12'hD51: soft_out = 32'h0000B6BB; // x = -10.7344, f(x) = 0.0000
    12'hD52: soft_out = 32'h0000B99C; // x = -10.7188, f(x) = 0.0000
    12'hD53: soft_out = 32'h0000BC88; // x = -10.7031, f(x) = 0.0000
    12'hD54: soft_out = 32'h0000BF80; // x = -10.6875, f(x) = 0.0000
    12'hD55: soft_out = 32'h0000C284; // x = -10.6719, f(x) = 0.0000
    12'hD56: soft_out = 32'h0000C594; // x = -10.6562, f(x) = 0.0000
    12'hD57: soft_out = 32'h0000C8B1; // x = -10.6406, f(x) = 0.0000
    12'hD58: soft_out = 32'h0000CBDA; // x = -10.6250, f(x) = 0.0000
    12'hD59: soft_out = 32'h0000CF0F; // x = -10.6094, f(x) = 0.0000
    12'hD5A: soft_out = 32'h0000D252; // x = -10.5938, f(x) = 0.0000
    12'hD5B: soft_out = 32'h0000D5A2; // x = -10.5781, f(x) = 0.0000
    12'hD5C: soft_out = 32'h0000D8FF; // x = -10.5625, f(x) = 0.0000
    12'hD5D: soft_out = 32'h0000DC6A; // x = -10.5469, f(x) = 0.0000
    12'hD5E: soft_out = 32'h0000DFE3; // x = -10.5312, f(x) = 0.0000
    12'hD5F: soft_out = 32'h0000E369; // x = -10.5156, f(x) = 0.0000
    12'hD60: soft_out = 32'h0000E6FE; // x = -10.5000, f(x) = 0.0000
    12'hD61: soft_out = 32'h0000EAA1; // x = -10.4844, f(x) = 0.0000
    12'hD62: soft_out = 32'h0000EE53; // x = -10.4688, f(x) = 0.0000
    12'hD63: soft_out = 32'h0000F214; // x = -10.4531, f(x) = 0.0000
    12'hD64: soft_out = 32'h0000F5E4; // x = -10.4375, f(x) = 0.0000
    12'hD65: soft_out = 32'h0000F9C3; // x = -10.4219, f(x) = 0.0000
    12'hD66: soft_out = 32'h0000FDB2; // x = -10.4062, f(x) = 0.0000
    12'hD67: soft_out = 32'h000101B1; // x = -10.3906, f(x) = 0.0000
    12'hD68: soft_out = 32'h000105C0; // x = -10.3750, f(x) = 0.0000
    12'hD69: soft_out = 32'h000109DF; // x = -10.3594, f(x) = 0.0000
    12'hD6A: soft_out = 32'h00010E0F; // x = -10.3438, f(x) = 0.0000
    12'hD6B: soft_out = 32'h0001124F; // x = -10.3281, f(x) = 0.0000
    12'hD6C: soft_out = 32'h000116A1; // x = -10.3125, f(x) = 0.0000
    12'hD6D: soft_out = 32'h00011B05; // x = -10.2969, f(x) = 0.0000
    12'hD6E: soft_out = 32'h00011F7A; // x = -10.2812, f(x) = 0.0000
    12'hD6F: soft_out = 32'h00012400; // x = -10.2656, f(x) = 0.0000
    12'hD70: soft_out = 32'h0001289A; // x = -10.2500, f(x) = 0.0000
    12'hD71: soft_out = 32'h00012D45; // x = -10.2344, f(x) = 0.0000
    12'hD72: soft_out = 32'h00013204; // x = -10.2188, f(x) = 0.0000
    12'hD73: soft_out = 32'h000136D6; // x = -10.2031, f(x) = 0.0000
    12'hD74: soft_out = 32'h00013BBB; // x = -10.1875, f(x) = 0.0000
    12'hD75: soft_out = 32'h000140B4; // x = -10.1719, f(x) = 0.0000
    12'hD76: soft_out = 32'h000145C0; // x = -10.1562, f(x) = 0.0000
    12'hD77: soft_out = 32'h00014AE2; // x = -10.1406, f(x) = 0.0000
    12'hD78: soft_out = 32'h00015018; // x = -10.1250, f(x) = 0.0000
    12'hD79: soft_out = 32'h00015562; // x = -10.1094, f(x) = 0.0000
    12'hD7A: soft_out = 32'h00015AC3; // x = -10.0938, f(x) = 0.0000
    12'hD7B: soft_out = 32'h00016039; // x = -10.0781, f(x) = 0.0000
    12'hD7C: soft_out = 32'h000165C5; // x = -10.0625, f(x) = 0.0000
    12'hD7D: soft_out = 32'h00016B67; // x = -10.0469, f(x) = 0.0000
    12'hD7E: soft_out = 32'h00017120; // x = -10.0312, f(x) = 0.0000
    12'hD7F: soft_out = 32'h000176F0; // x = -10.0156, f(x) = 0.0000
    12'hD80: soft_out = 32'h00017CD8; // x = -10.0000, f(x) = 0.0000
    12'hD81: soft_out = 32'h000182D7; // x = -9.9844, f(x) = 0.0000
    12'hD82: soft_out = 32'h000188EE; // x = -9.9688, f(x) = 0.0000
    12'hD83: soft_out = 32'h00018F1F; // x = -9.9531, f(x) = 0.0000
    12'hD84: soft_out = 32'h00019568; // x = -9.9375, f(x) = 0.0000
    12'hD85: soft_out = 32'h00019BCA; // x = -9.9219, f(x) = 0.0000
    12'hD86: soft_out = 32'h0001A246; // x = -9.9062, f(x) = 0.0000
    12'hD87: soft_out = 32'h0001A8DC; // x = -9.8906, f(x) = 0.0001
    12'hD88: soft_out = 32'h0001AF8D; // x = -9.8750, f(x) = 0.0001
    12'hD89: soft_out = 32'h0001B659; // x = -9.8594, f(x) = 0.0001
    12'hD8A: soft_out = 32'h0001BD40; // x = -9.8438, f(x) = 0.0001
    12'hD8B: soft_out = 32'h0001C443; // x = -9.8281, f(x) = 0.0001
    12'hD8C: soft_out = 32'h0001CB62; // x = -9.8125, f(x) = 0.0001
    12'hD8D: soft_out = 32'h0001D29E; // x = -9.7969, f(x) = 0.0001
    12'hD8E: soft_out = 32'h0001D9F7; // x = -9.7812, f(x) = 0.0001
    12'hD8F: soft_out = 32'h0001E16E; // x = -9.7656, f(x) = 0.0001
    12'hD90: soft_out = 32'h0001E903; // x = -9.7500, f(x) = 0.0001
    12'hD91: soft_out = 32'h0001F0B6; // x = -9.7344, f(x) = 0.0001
    12'hD92: soft_out = 32'h0001F889; // x = -9.7188, f(x) = 0.0001
    12'hD93: soft_out = 32'h0002007B; // x = -9.7031, f(x) = 0.0001
    12'hD94: soft_out = 32'h0002088D; // x = -9.6875, f(x) = 0.0001
    12'hD95: soft_out = 32'h000210BF; // x = -9.6719, f(x) = 0.0001
    12'hD96: soft_out = 32'h00021913; // x = -9.6562, f(x) = 0.0001
    12'hD97: soft_out = 32'h00022188; // x = -9.6406, f(x) = 0.0001
    12'hD98: soft_out = 32'h00022A1F; // x = -9.6250, f(x) = 0.0001
    12'hD99: soft_out = 32'h000232D9; // x = -9.6094, f(x) = 0.0001
    12'hD9A: soft_out = 32'h00023BB6; // x = -9.5938, f(x) = 0.0001
    12'hD9B: soft_out = 32'h000244B7; // x = -9.5781, f(x) = 0.0001
    12'hD9C: soft_out = 32'h00024DDC; // x = -9.5625, f(x) = 0.0001
    12'hD9D: soft_out = 32'h00025726; // x = -9.5469, f(x) = 0.0001
    12'hD9E: soft_out = 32'h00026096; // x = -9.5312, f(x) = 0.0001
    12'hD9F: soft_out = 32'h00026A2B; // x = -9.5156, f(x) = 0.0001
    12'hDA0: soft_out = 32'h000273E7; // x = -9.5000, f(x) = 0.0001
    12'hDA1: soft_out = 32'h00027DCA; // x = -9.4844, f(x) = 0.0001
    12'hDA2: soft_out = 32'h000287D6; // x = -9.4688, f(x) = 0.0001
    12'hDA3: soft_out = 32'h00029209; // x = -9.4531, f(x) = 0.0001
    12'hDA4: soft_out = 32'h00029C66; // x = -9.4375, f(x) = 0.0001
    12'hDA5: soft_out = 32'h0002A6ED; // x = -9.4219, f(x) = 0.0001
    12'hDA6: soft_out = 32'h0002B19E; // x = -9.4062, f(x) = 0.0001
    12'hDA7: soft_out = 32'h0002BC7A; // x = -9.3906, f(x) = 0.0001
    12'hDA8: soft_out = 32'h0002C782; // x = -9.3750, f(x) = 0.0001
    12'hDA9: soft_out = 32'h0002D2B6; // x = -9.3594, f(x) = 0.0001
    12'hDAA: soft_out = 32'h0002DE18; // x = -9.3438, f(x) = 0.0001
    12'hDAB: soft_out = 32'h0002E9A7; // x = -9.3281, f(x) = 0.0001
    12'hDAC: soft_out = 32'h0002F565; // x = -9.3125, f(x) = 0.0001
    12'hDAD: soft_out = 32'h00030153; // x = -9.2969, f(x) = 0.0001
    12'hDAE: soft_out = 32'h00030D70; // x = -9.2812, f(x) = 0.0001
    12'hDAF: soft_out = 32'h000319BE; // x = -9.2656, f(x) = 0.0001
    12'hDB0: soft_out = 32'h0003263E; // x = -9.2500, f(x) = 0.0001
    12'hDB1: soft_out = 32'h000332F0; // x = -9.2344, f(x) = 0.0001
    12'hDB2: soft_out = 32'h00033FD6; // x = -9.2188, f(x) = 0.0001
    12'hDB3: soft_out = 32'h00034CEF; // x = -9.2031, f(x) = 0.0001
    12'hDB4: soft_out = 32'h00035A3E; // x = -9.1875, f(x) = 0.0001
    12'hDB5: soft_out = 32'h000367C2; // x = -9.1719, f(x) = 0.0001
    12'hDB6: soft_out = 32'h0003757C; // x = -9.1562, f(x) = 0.0001
    12'hDB7: soft_out = 32'h0003836E; // x = -9.1406, f(x) = 0.0001
    12'hDB8: soft_out = 32'h00039198; // x = -9.1250, f(x) = 0.0001
    12'hDB9: soft_out = 32'h00039FFB; // x = -9.1094, f(x) = 0.0001
    12'hDBA: soft_out = 32'h0003AE98; // x = -9.0938, f(x) = 0.0001
    12'hDBB: soft_out = 32'h0003BD70; // x = -9.0781, f(x) = 0.0001
    12'hDBC: soft_out = 32'h0003CC84; // x = -9.0625, f(x) = 0.0001
    12'hDBD: soft_out = 32'h0003DBD4; // x = -9.0469, f(x) = 0.0001
    12'hDBE: soft_out = 32'h0003EB63; // x = -9.0312, f(x) = 0.0001
    12'hDBF: soft_out = 32'h0003FB30; // x = -9.0156, f(x) = 0.0001
    12'hDC0: soft_out = 32'h00040B3D; // x = -9.0000, f(x) = 0.0001
    12'hDC1: soft_out = 32'h00041B8A; // x = -8.9844, f(x) = 0.0001
    12'hDC2: soft_out = 32'h00042C19; // x = -8.9688, f(x) = 0.0001
    12'hDC3: soft_out = 32'h00043CEB; // x = -8.9531, f(x) = 0.0001
    12'hDC4: soft_out = 32'h00044E01; // x = -8.9375, f(x) = 0.0001
    12'hDC5: soft_out = 32'h00045F5C; // x = -8.9219, f(x) = 0.0001
    12'hDC6: soft_out = 32'h000470FC; // x = -8.9062, f(x) = 0.0001
    12'hDC7: soft_out = 32'h000482E4; // x = -8.8906, f(x) = 0.0001
    12'hDC8: soft_out = 32'h00049514; // x = -8.8750, f(x) = 0.0001
    12'hDC9: soft_out = 32'h0004A78D; // x = -8.8594, f(x) = 0.0001
    12'hDCA: soft_out = 32'h0004BA50; // x = -8.8438, f(x) = 0.0001
    12'hDCB: soft_out = 32'h0004CD60; // x = -8.8281, f(x) = 0.0001
    12'hDCC: soft_out = 32'h0004E0BC; // x = -8.8125, f(x) = 0.0001
    12'hDCD: soft_out = 32'h0004F466; // x = -8.7969, f(x) = 0.0002
    12'hDCE: soft_out = 32'h0005085F; // x = -8.7812, f(x) = 0.0002
    12'hDCF: soft_out = 32'h00051CA9; // x = -8.7656, f(x) = 0.0002
    12'hDD0: soft_out = 32'h00053145; // x = -8.7500, f(x) = 0.0002
    12'hDD1: soft_out = 32'h00054634; // x = -8.7344, f(x) = 0.0002
    12'hDD2: soft_out = 32'h00055B77; // x = -8.7188, f(x) = 0.0002
    12'hDD3: soft_out = 32'h00057110; // x = -8.7031, f(x) = 0.0002
    12'hDD4: soft_out = 32'h00058700; // x = -8.6875, f(x) = 0.0002
    12'hDD5: soft_out = 32'h00059D49; // x = -8.6719, f(x) = 0.0002
    12'hDD6: soft_out = 32'h0005B3EB; // x = -8.6562, f(x) = 0.0002
    12'hDD7: soft_out = 32'h0005CAE8; // x = -8.6406, f(x) = 0.0002
    12'hDD8: soft_out = 32'h0005E243; // x = -8.6250, f(x) = 0.0002
    12'hDD9: soft_out = 32'h0005F9FB; // x = -8.6094, f(x) = 0.0002
    12'hDDA: soft_out = 32'h00061213; // x = -8.5938, f(x) = 0.0002
    12'hDDB: soft_out = 32'h00062A8C; // x = -8.5781, f(x) = 0.0002
    12'hDDC: soft_out = 32'h00064368; // x = -8.5625, f(x) = 0.0002
    12'hDDD: soft_out = 32'h00065CA8; // x = -8.5469, f(x) = 0.0002
    12'hDDE: soft_out = 32'h0006764E; // x = -8.5312, f(x) = 0.0002
    12'hDDF: soft_out = 32'h0006905B; // x = -8.5156, f(x) = 0.0002
    12'hDE0: soft_out = 32'h0006AAD1; // x = -8.5000, f(x) = 0.0002
    12'hDE1: soft_out = 32'h0006C5B2; // x = -8.4844, f(x) = 0.0002
    12'hDE2: soft_out = 32'h0006E0FF; // x = -8.4688, f(x) = 0.0002
    12'hDE3: soft_out = 32'h0006FCBA; // x = -8.4531, f(x) = 0.0002
    12'hDE4: soft_out = 32'h000718E6; // x = -8.4375, f(x) = 0.0002
    12'hDE5: soft_out = 32'h00073582; // x = -8.4219, f(x) = 0.0002
    12'hDE6: soft_out = 32'h00075292; // x = -8.4062, f(x) = 0.0002
    12'hDE7: soft_out = 32'h00077017; // x = -8.3906, f(x) = 0.0002
    12'hDE8: soft_out = 32'h00078E14; // x = -8.3750, f(x) = 0.0002
    12'hDE9: soft_out = 32'h0007AC89; // x = -8.3594, f(x) = 0.0002
    12'hDEA: soft_out = 32'h0007CB78; // x = -8.3438, f(x) = 0.0002
    12'hDEB: soft_out = 32'h0007EAE5; // x = -8.3281, f(x) = 0.0002
    12'hDEC: soft_out = 32'h00080AD0; // x = -8.3125, f(x) = 0.0002
    12'hDED: soft_out = 32'h00082B3C; // x = -8.2969, f(x) = 0.0002
    12'hDEE: soft_out = 32'h00084C2B; // x = -8.2812, f(x) = 0.0003
    12'hDEF: soft_out = 32'h00086D9E; // x = -8.2656, f(x) = 0.0003
    12'hDF0: soft_out = 32'h00088F98; // x = -8.2500, f(x) = 0.0003
    12'hDF1: soft_out = 32'h0008B21C; // x = -8.2344, f(x) = 0.0003
    12'hDF2: soft_out = 32'h0008D52A; // x = -8.2188, f(x) = 0.0003
    12'hDF3: soft_out = 32'h0008F8C6; // x = -8.2031, f(x) = 0.0003
    12'hDF4: soft_out = 32'h00091CF1; // x = -8.1875, f(x) = 0.0003
    12'hDF5: soft_out = 32'h000941AE; // x = -8.1719, f(x) = 0.0003
    12'hDF6: soft_out = 32'h000966FF; // x = -8.1562, f(x) = 0.0003
    12'hDF7: soft_out = 32'h00098CE7; // x = -8.1406, f(x) = 0.0003
    12'hDF8: soft_out = 32'h0009B367; // x = -8.1250, f(x) = 0.0003
    12'hDF9: soft_out = 32'h0009DA83; // x = -8.1094, f(x) = 0.0003
    12'hDFA: soft_out = 32'h000A023C; // x = -8.0938, f(x) = 0.0003
    12'hDFB: soft_out = 32'h000A2A96; // x = -8.0781, f(x) = 0.0003
    12'hDFC: soft_out = 32'h000A5392; // x = -8.0625, f(x) = 0.0003
    12'hDFD: soft_out = 32'h000A7D33; // x = -8.0469, f(x) = 0.0003
    12'hDFE: soft_out = 32'h000AA77C; // x = -8.0312, f(x) = 0.0003
    12'hDFF: soft_out = 32'h000AD270; // x = -8.0156, f(x) = 0.0003
    12'hE00: soft_out = 32'h000AFE11; // x = -8.0000, f(x) = 0.0003
    12'hE01: soft_out = 32'h000B2A61; // x = -7.9844, f(x) = 0.0003
    12'hE02: soft_out = 32'h000B5764; // x = -7.9688, f(x) = 0.0003
    12'hE03: soft_out = 32'h000B851D; // x = -7.9531, f(x) = 0.0004
    12'hE04: soft_out = 32'h000BB38E; // x = -7.9375, f(x) = 0.0004
    12'hE05: soft_out = 32'h000BE2BB; // x = -7.9219, f(x) = 0.0004
    12'hE06: soft_out = 32'h000C12A5; // x = -7.9062, f(x) = 0.0004
    12'hE07: soft_out = 32'h000C4351; // x = -7.8906, f(x) = 0.0004
    12'hE08: soft_out = 32'h000C74C1; // x = -7.8750, f(x) = 0.0004
    12'hE09: soft_out = 32'h000CA6F8; // x = -7.8594, f(x) = 0.0004
    12'hE0A: soft_out = 32'h000CD9FA; // x = -7.8438, f(x) = 0.0004
    12'hE0B: soft_out = 32'h000D0DC9; // x = -7.8281, f(x) = 0.0004
    12'hE0C: soft_out = 32'h000D4269; // x = -7.8125, f(x) = 0.0004
    12'hE0D: soft_out = 32'h000D77DD; // x = -7.7969, f(x) = 0.0004
    12'hE0E: soft_out = 32'h000DAE29; // x = -7.7812, f(x) = 0.0004
    12'hE0F: soft_out = 32'h000DE550; // x = -7.7656, f(x) = 0.0004
    12'hE10: soft_out = 32'h000E1D55; // x = -7.7500, f(x) = 0.0004
    12'hE11: soft_out = 32'h000E563B; // x = -7.7344, f(x) = 0.0004
    12'hE12: soft_out = 32'h000E9008; // x = -7.7188, f(x) = 0.0004
    12'hE13: soft_out = 32'h000ECABD; // x = -7.7031, f(x) = 0.0005
    12'hE14: soft_out = 32'h000F065F; // x = -7.6875, f(x) = 0.0005
    12'hE15: soft_out = 32'h000F42F1; // x = -7.6719, f(x) = 0.0005
    12'hE16: soft_out = 32'h000F8078; // x = -7.6562, f(x) = 0.0005
    12'hE17: soft_out = 32'h000FBEF6; // x = -7.6406, f(x) = 0.0005
    12'hE18: soft_out = 32'h000FFE71; // x = -7.6250, f(x) = 0.0005
    12'hE19: soft_out = 32'h00103EEB; // x = -7.6094, f(x) = 0.0005
    12'hE1A: soft_out = 32'h00108069; // x = -7.5938, f(x) = 0.0005
    12'hE1B: soft_out = 32'h0010C2F0; // x = -7.5781, f(x) = 0.0005
    12'hE1C: soft_out = 32'h00110682; // x = -7.5625, f(x) = 0.0005
    12'hE1D: soft_out = 32'h00114B25; // x = -7.5469, f(x) = 0.0005
    12'hE1E: soft_out = 32'h001190DD; // x = -7.5312, f(x) = 0.0005
    12'hE1F: soft_out = 32'h0011D7AD; // x = -7.5156, f(x) = 0.0005
    12'hE20: soft_out = 32'h00121F9C; // x = -7.5000, f(x) = 0.0006
    12'hE21: soft_out = 32'h001268AC; // x = -7.4844, f(x) = 0.0006
    12'hE22: soft_out = 32'h0012B2E3; // x = -7.4688, f(x) = 0.0006
    12'hE23: soft_out = 32'h0012FE44; // x = -7.4531, f(x) = 0.0006
    12'hE24: soft_out = 32'h00134AD6; // x = -7.4375, f(x) = 0.0006
    12'hE25: soft_out = 32'h0013989D; // x = -7.4219, f(x) = 0.0006
    12'hE26: soft_out = 32'h0013E79D; // x = -7.4062, f(x) = 0.0006
    12'hE27: soft_out = 32'h001437DB; // x = -7.3906, f(x) = 0.0006
    12'hE28: soft_out = 32'h0014895D; // x = -7.3750, f(x) = 0.0006
    12'hE29: soft_out = 32'h0014DC28; // x = -7.3594, f(x) = 0.0006
    12'hE2A: soft_out = 32'h00153040; // x = -7.3438, f(x) = 0.0006
    12'hE2B: soft_out = 32'h001585AC; // x = -7.3281, f(x) = 0.0007
    12'hE2C: soft_out = 32'h0015DC6F; // x = -7.3125, f(x) = 0.0007
    12'hE2D: soft_out = 32'h00163491; // x = -7.2969, f(x) = 0.0007
    12'hE2E: soft_out = 32'h00168E16; // x = -7.2812, f(x) = 0.0007
    12'hE2F: soft_out = 32'h0016E904; // x = -7.2656, f(x) = 0.0007
    12'hE30: soft_out = 32'h00174560; // x = -7.2500, f(x) = 0.0007
    12'hE31: soft_out = 32'h0017A331; // x = -7.2344, f(x) = 0.0007
    12'hE32: soft_out = 32'h0018027B; // x = -7.2188, f(x) = 0.0007
    12'hE33: soft_out = 32'h00186346; // x = -7.2031, f(x) = 0.0007
    12'hE34: soft_out = 32'h0018C598; // x = -7.1875, f(x) = 0.0008
    12'hE35: soft_out = 32'h00192975; // x = -7.1719, f(x) = 0.0008
    12'hE36: soft_out = 32'h00198EE5; // x = -7.1562, f(x) = 0.0008
    12'hE37: soft_out = 32'h0019F5EE; // x = -7.1406, f(x) = 0.0008
    12'hE38: soft_out = 32'h001A5E97; // x = -7.1250, f(x) = 0.0008
    12'hE39: soft_out = 32'h001AC8E5; // x = -7.1094, f(x) = 0.0008
    12'hE3A: soft_out = 32'h001B34E0; // x = -7.0938, f(x) = 0.0008
    12'hE3B: soft_out = 32'h001BA28F; // x = -7.0781, f(x) = 0.0008
    12'hE3C: soft_out = 32'h001C11F7; // x = -7.0625, f(x) = 0.0009
    12'hE3D: soft_out = 32'h001C8321; // x = -7.0469, f(x) = 0.0009
    12'hE3E: soft_out = 32'h001CF613; // x = -7.0312, f(x) = 0.0009
    12'hE3F: soft_out = 32'h001D6AD4; // x = -7.0156, f(x) = 0.0009
    12'hE40: soft_out = 32'h001DE16C; // x = -7.0000, f(x) = 0.0009
    12'hE41: soft_out = 32'h001E59E2; // x = -6.9844, f(x) = 0.0009
    12'hE42: soft_out = 32'h001ED43D; // x = -6.9688, f(x) = 0.0009
    12'hE43: soft_out = 32'h001F5086; // x = -6.9531, f(x) = 0.0010
    12'hE44: soft_out = 32'h001FCEC4; // x = -6.9375, f(x) = 0.0010
    12'hE45: soft_out = 32'h00204EFF; // x = -6.9219, f(x) = 0.0010
    12'hE46: soft_out = 32'h0020D13F; // x = -6.9062, f(x) = 0.0010
    12'hE47: soft_out = 32'h0021558C; // x = -6.8906, f(x) = 0.0010
    12'hE48: soft_out = 32'h0021DBEE; // x = -6.8750, f(x) = 0.0010
    12'hE49: soft_out = 32'h0022646E; // x = -6.8594, f(x) = 0.0010
    12'hE4A: soft_out = 32'h0022EF14; // x = -6.8438, f(x) = 0.0011
    12'hE4B: soft_out = 32'h00237BE9; // x = -6.8281, f(x) = 0.0011
    12'hE4C: soft_out = 32'h00240AF6; // x = -6.8125, f(x) = 0.0011
    12'hE4D: soft_out = 32'h00249C44; // x = -6.7969, f(x) = 0.0011
    12'hE4E: soft_out = 32'h00252FDC; // x = -6.7812, f(x) = 0.0011
    12'hE4F: soft_out = 32'h0025C5C6; // x = -6.7656, f(x) = 0.0012
    12'hE50: soft_out = 32'h00265E0D; // x = -6.7500, f(x) = 0.0012
    12'hE51: soft_out = 32'h0026F8BA; // x = -6.7344, f(x) = 0.0012
    12'hE52: soft_out = 32'h002795D6; // x = -6.7188, f(x) = 0.0012
    12'hE53: soft_out = 32'h0028356C; // x = -6.7031, f(x) = 0.0012
    12'hE54: soft_out = 32'h0028D785; // x = -6.6875, f(x) = 0.0012
    12'hE55: soft_out = 32'h00297C2B; // x = -6.6719, f(x) = 0.0013
    12'hE56: soft_out = 32'h002A2369; // x = -6.6562, f(x) = 0.0013
    12'hE57: soft_out = 32'h002ACD4A; // x = -6.6406, f(x) = 0.0013
    12'hE58: soft_out = 32'h002B79D7; // x = -6.6250, f(x) = 0.0013
    12'hE59: soft_out = 32'h002C291C; // x = -6.6094, f(x) = 0.0013
    12'hE5A: soft_out = 32'h002CDB24; // x = -6.5938, f(x) = 0.0014
    12'hE5B: soft_out = 32'h002D8FF9; // x = -6.5781, f(x) = 0.0014
    12'hE5C: soft_out = 32'h002E47A7; // x = -6.5625, f(x) = 0.0014
    12'hE5D: soft_out = 32'h002F023A; // x = -6.5469, f(x) = 0.0014
    12'hE5E: soft_out = 32'h002FBFBD; // x = -6.5312, f(x) = 0.0015
    12'hE5F: soft_out = 32'h0030803C; // x = -6.5156, f(x) = 0.0015
    12'hE60: soft_out = 32'h003143C3; // x = -6.5000, f(x) = 0.0015
    12'hE61: soft_out = 32'h00320A5E; // x = -6.4844, f(x) = 0.0015
    12'hE62: soft_out = 32'h0032D41A; // x = -6.4688, f(x) = 0.0016
    12'hE63: soft_out = 32'h0033A103; // x = -6.4531, f(x) = 0.0016
    12'hE64: soft_out = 32'h00347127; // x = -6.4375, f(x) = 0.0016
    12'hE65: soft_out = 32'h00354491; // x = -6.4219, f(x) = 0.0016
    12'hE66: soft_out = 32'h00361B50; // x = -6.4062, f(x) = 0.0017
    12'hE67: soft_out = 32'h0036F570; // x = -6.3906, f(x) = 0.0017
    12'hE68: soft_out = 32'h0037D300; // x = -6.3750, f(x) = 0.0017
    12'hE69: soft_out = 32'h0038B40D; // x = -6.3594, f(x) = 0.0017
    12'hE6A: soft_out = 32'h003998A5; // x = -6.3438, f(x) = 0.0018
    12'hE6B: soft_out = 32'h003A80D7; // x = -6.3281, f(x) = 0.0018
    12'hE6C: soft_out = 32'h003B6CB0; // x = -6.3125, f(x) = 0.0018
    12'hE6D: soft_out = 32'h003C5C41; // x = -6.2969, f(x) = 0.0018
    12'hE6E: soft_out = 32'h003D4F97; // x = -6.2812, f(x) = 0.0019
    12'hE6F: soft_out = 32'h003E46C3; // x = -6.2656, f(x) = 0.0019
    12'hE70: soft_out = 32'h003F41D3; // x = -6.2500, f(x) = 0.0019
    12'hE71: soft_out = 32'h004040D7; // x = -6.2344, f(x) = 0.0020
    12'hE72: soft_out = 32'h004143DF; // x = -6.2188, f(x) = 0.0020
    12'hE73: soft_out = 32'h00424AFB; // x = -6.2031, f(x) = 0.0020
    12'hE74: soft_out = 32'h0043563C; // x = -6.1875, f(x) = 0.0021
    12'hE75: soft_out = 32'h004465B3; // x = -6.1719, f(x) = 0.0021
    12'hE76: soft_out = 32'h0045796F; // x = -6.1562, f(x) = 0.0021
    12'hE77: soft_out = 32'h00469184; // x = -6.1406, f(x) = 0.0022
    12'hE78: soft_out = 32'h0047AE01; // x = -6.1250, f(x) = 0.0022
    12'hE79: soft_out = 32'h0048CEFA; // x = -6.1094, f(x) = 0.0022
    12'hE7A: soft_out = 32'h0049F47F; // x = -6.0938, f(x) = 0.0023
    12'hE7B: soft_out = 32'h004B1EA4; // x = -6.0781, f(x) = 0.0023
    12'hE7C: soft_out = 32'h004C4D7B; // x = -6.0625, f(x) = 0.0023
    12'hE7D: soft_out = 32'h004D8116; // x = -6.0469, f(x) = 0.0024
    12'hE7E: soft_out = 32'h004EB98A; // x = -6.0312, f(x) = 0.0024
    12'hE7F: soft_out = 32'h004FF6E9; // x = -6.0156, f(x) = 0.0024
    12'hE80: soft_out = 32'h00513948; // x = -6.0000, f(x) = 0.0025
    12'hE81: soft_out = 32'h005280BA; // x = -5.9844, f(x) = 0.0025
    12'hE82: soft_out = 32'h0053CD54; // x = -5.9688, f(x) = 0.0026
    12'hE83: soft_out = 32'h00551F2C; // x = -5.9531, f(x) = 0.0026
    12'hE84: soft_out = 32'h00567655; // x = -5.9375, f(x) = 0.0026
    12'hE85: soft_out = 32'h0057D2E6; // x = -5.9219, f(x) = 0.0027
    12'hE86: soft_out = 32'h005934F3; // x = -5.9062, f(x) = 0.0027
    12'hE87: soft_out = 32'h005A9C95; // x = -5.8906, f(x) = 0.0028
    12'hE88: soft_out = 32'h005C09E0; // x = -5.8750, f(x) = 0.0028
    12'hE89: soft_out = 32'h005D7CEB; // x = -5.8594, f(x) = 0.0029
    12'hE8A: soft_out = 32'h005EF5CF; // x = -5.8438, f(x) = 0.0029
    12'hE8B: soft_out = 32'h006074A2; // x = -5.8281, f(x) = 0.0029
    12'hE8C: soft_out = 32'h0061F97C; // x = -5.8125, f(x) = 0.0030
    12'hE8D: soft_out = 32'h00638476; // x = -5.7969, f(x) = 0.0030
    12'hE8E: soft_out = 32'h006515A8; // x = -5.7812, f(x) = 0.0031
    12'hE8F: soft_out = 32'h0066AD2B; // x = -5.7656, f(x) = 0.0031
    12'hE90: soft_out = 32'h00684B1A; // x = -5.7500, f(x) = 0.0032
    12'hE91: soft_out = 32'h0069EF8D; // x = -5.7344, f(x) = 0.0032
    12'hE92: soft_out = 32'h006B9A9F; // x = -5.7188, f(x) = 0.0033
    12'hE93: soft_out = 32'h006D4C6B; // x = -5.7031, f(x) = 0.0033
    12'hE94: soft_out = 32'h006F050B; // x = -5.6875, f(x) = 0.0034
    12'hE95: soft_out = 32'h0070C49C; // x = -5.6719, f(x) = 0.0034
    12'hE96: soft_out = 32'h00728B3A; // x = -5.6562, f(x) = 0.0035
    12'hE97: soft_out = 32'h00745900; // x = -5.6406, f(x) = 0.0036
    12'hE98: soft_out = 32'h00762E0B; // x = -5.6250, f(x) = 0.0036
    12'hE99: soft_out = 32'h00780A7A; // x = -5.6094, f(x) = 0.0037
    12'hE9A: soft_out = 32'h0079EE69; // x = -5.5938, f(x) = 0.0037
    12'hE9B: soft_out = 32'h007BD9F7; // x = -5.5781, f(x) = 0.0038
    12'hE9C: soft_out = 32'h007DCD43; // x = -5.5625, f(x) = 0.0038
    12'hE9D: soft_out = 32'h007FC86C; // x = -5.5469, f(x) = 0.0039
    12'hE9E: soft_out = 32'h0081CB91; // x = -5.5312, f(x) = 0.0040
    12'hE9F: soft_out = 32'h0083D6D3; // x = -5.5156, f(x) = 0.0040
    12'hEA0: soft_out = 32'h0085EA53; // x = -5.5000, f(x) = 0.0041
    12'hEA1: soft_out = 32'h00880631; // x = -5.4844, f(x) = 0.0042
    12'hEA2: soft_out = 32'h008A2A90; // x = -5.4688, f(x) = 0.0042
    12'hEA3: soft_out = 32'h008C5791; // x = -5.4531, f(x) = 0.0043
    12'hEA4: soft_out = 32'h008E8D58; // x = -5.4375, f(x) = 0.0044
    12'hEA5: soft_out = 32'h0090CC08; // x = -5.4219, f(x) = 0.0044
    12'hEA6: soft_out = 32'h009313C4; // x = -5.4062, f(x) = 0.0045
    12'hEA7: soft_out = 32'h009564B2; // x = -5.3906, f(x) = 0.0046
    12'hEA8: soft_out = 32'h0097BEF6; // x = -5.3750, f(x) = 0.0046
    12'hEA9: soft_out = 32'h009A22B6; // x = -5.3594, f(x) = 0.0047
    12'hEAA: soft_out = 32'h009C9019; // x = -5.3438, f(x) = 0.0048
    12'hEAB: soft_out = 32'h009F0744; // x = -5.3281, f(x) = 0.0049
    12'hEAC: soft_out = 32'h00A18860; // x = -5.3125, f(x) = 0.0049
    12'hEAD: soft_out = 32'h00A41395; // x = -5.2969, f(x) = 0.0050
    12'hEAE: soft_out = 32'h00A6A90B; // x = -5.2812, f(x) = 0.0051
    12'hEAF: soft_out = 32'h00A948EB; // x = -5.2656, f(x) = 0.0052
    12'hEB0: soft_out = 32'h00ABF360; // x = -5.2500, f(x) = 0.0052
    12'hEB1: soft_out = 32'h00AEA894; // x = -5.2344, f(x) = 0.0053
    12'hEB2: soft_out = 32'h00B168B3; // x = -5.2188, f(x) = 0.0054
    12'hEB3: soft_out = 32'h00B433E9; // x = -5.2031, f(x) = 0.0055
    12'hEB4: soft_out = 32'h00B70A61; // x = -5.1875, f(x) = 0.0056
    12'hEB5: soft_out = 32'h00B9EC4B; // x = -5.1719, f(x) = 0.0057
    12'hEB6: soft_out = 32'h00BCD9D3; // x = -5.1562, f(x) = 0.0058
    12'hEB7: soft_out = 32'h00BFD329; // x = -5.1406, f(x) = 0.0059
    12'hEB8: soft_out = 32'h00C2D87D; // x = -5.1250, f(x) = 0.0059
    12'hEB9: soft_out = 32'h00C5E9FD; // x = -5.1094, f(x) = 0.0060
    12'hEBA: soft_out = 32'h00C907DD; // x = -5.0938, f(x) = 0.0061
    12'hEBB: soft_out = 32'h00CC324D; // x = -5.0781, f(x) = 0.0062
    12'hEBC: soft_out = 32'h00CF6980; // x = -5.0625, f(x) = 0.0063
    12'hEBD: soft_out = 32'h00D2ADAA; // x = -5.0469, f(x) = 0.0064
    12'hEBE: soft_out = 32'h00D5FEFF; // x = -5.0312, f(x) = 0.0065
    12'hEBF: soft_out = 32'h00D95DB4; // x = -5.0156, f(x) = 0.0066
    12'hEC0: soft_out = 32'h00DCC9FF; // x = -5.0000, f(x) = 0.0067
    12'hEC1: soft_out = 32'h00E04417; // x = -4.9844, f(x) = 0.0068
    12'hEC2: soft_out = 32'h00E3CC32; // x = -4.9688, f(x) = 0.0070
    12'hEC3: soft_out = 32'h00E7628B; // x = -4.9531, f(x) = 0.0071
    12'hEC4: soft_out = 32'h00EB075A; // x = -4.9375, f(x) = 0.0072
    12'hEC5: soft_out = 32'h00EEBAD9; // x = -4.9219, f(x) = 0.0073
    12'hEC6: soft_out = 32'h00F27D45; // x = -4.9062, f(x) = 0.0074
    12'hEC7: soft_out = 32'h00F64ED8; // x = -4.8906, f(x) = 0.0075
    12'hEC8: soft_out = 32'h00FA2FD0; // x = -4.8750, f(x) = 0.0076
    12'hEC9: soft_out = 32'h00FE206B; // x = -4.8594, f(x) = 0.0078
    12'hECA: soft_out = 32'h010220E9; // x = -4.8438, f(x) = 0.0079
    12'hECB: soft_out = 32'h01063188; // x = -4.8281, f(x) = 0.0080
    12'hECC: soft_out = 32'h010A528B; // x = -4.8125, f(x) = 0.0081
    12'hECD: soft_out = 32'h010E8432; // x = -4.7969, f(x) = 0.0083
    12'hECE: soft_out = 32'h0112C6C3; // x = -4.7812, f(x) = 0.0084
    12'hECF: soft_out = 32'h01171A7F; // x = -4.7656, f(x) = 0.0085
    12'hED0: soft_out = 32'h011B7FAE; // x = -4.7500, f(x) = 0.0087
    12'hED1: soft_out = 32'h011FF695; // x = -4.7344, f(x) = 0.0088
    12'hED2: soft_out = 32'h01247F7B; // x = -4.7188, f(x) = 0.0089
    12'hED3: soft_out = 32'h01291AA9; // x = -4.7031, f(x) = 0.0091
    12'hED4: soft_out = 32'h012DC869; // x = -4.6875, f(x) = 0.0092
    12'hED5: soft_out = 32'h01328905; // x = -4.6719, f(x) = 0.0094
    12'hED6: soft_out = 32'h01375CCA; // x = -4.6562, f(x) = 0.0095
    12'hED7: soft_out = 32'h013C4405; // x = -4.6406, f(x) = 0.0097
    12'hED8: soft_out = 32'h01413F05; // x = -4.6250, f(x) = 0.0098
    12'hED9: soft_out = 32'h01464E18; // x = -4.6094, f(x) = 0.0100
    12'hEDA: soft_out = 32'h014B7191; // x = -4.5938, f(x) = 0.0101
    12'hEDB: soft_out = 32'h0150A9C1; // x = -4.5781, f(x) = 0.0103
    12'hEDC: soft_out = 32'h0155F6FB; // x = -4.5625, f(x) = 0.0104
    12'hEDD: soft_out = 32'h015B5995; // x = -4.5469, f(x) = 0.0106
    12'hEDE: soft_out = 32'h0160D1E5; // x = -4.5312, f(x) = 0.0108
    12'hEDF: soft_out = 32'h01666041; // x = -4.5156, f(x) = 0.0109
    12'hEE0: soft_out = 32'h016C0504; // x = -4.5000, f(x) = 0.0111
    12'hEE1: soft_out = 32'h0171C088; // x = -4.4844, f(x) = 0.0113
    12'hEE2: soft_out = 32'h01779327; // x = -4.4688, f(x) = 0.0115
    12'hEE3: soft_out = 32'h017D7D40; // x = -4.4531, f(x) = 0.0116
    12'hEE4: soft_out = 32'h01837F31; // x = -4.4375, f(x) = 0.0118
    12'hEE5: soft_out = 32'h0189995A; // x = -4.4219, f(x) = 0.0120
    12'hEE6: soft_out = 32'h018FCC1D; // x = -4.4062, f(x) = 0.0122
    12'hEE7: soft_out = 32'h019617DC; // x = -4.3906, f(x) = 0.0124
    12'hEE8: soft_out = 32'h019C7CFE; // x = -4.3750, f(x) = 0.0126
    12'hEE9: soft_out = 32'h01A2FBE7; // x = -4.3594, f(x) = 0.0128
    12'hEEA: soft_out = 32'h01A99500; // x = -4.3438, f(x) = 0.0130
    12'hEEB: soft_out = 32'h01B048B2; // x = -4.3281, f(x) = 0.0132
    12'hEEC: soft_out = 32'h01B71769; // x = -4.3125, f(x) = 0.0134
    12'hEED: soft_out = 32'h01BE0192; // x = -4.2969, f(x) = 0.0136
    12'hEEE: soft_out = 32'h01C5079B; // x = -4.2812, f(x) = 0.0138
    12'hEEF: soft_out = 32'h01CC29F5; // x = -4.2656, f(x) = 0.0140
    12'hEF0: soft_out = 32'h01D36911; // x = -4.2500, f(x) = 0.0143
    12'hEF1: soft_out = 32'h01DAC564; // x = -4.2344, f(x) = 0.0145
    12'hEF2: soft_out = 32'h01E23F64; // x = -4.2188, f(x) = 0.0147
    12'hEF3: soft_out = 32'h01E9D787; // x = -4.2031, f(x) = 0.0149
    12'hEF4: soft_out = 32'h01F18E49; // x = -4.1875, f(x) = 0.0152
    12'hEF5: soft_out = 32'h01F96423; // x = -4.1719, f(x) = 0.0154
    12'hEF6: soft_out = 32'h02015994; // x = -4.1562, f(x) = 0.0157
    12'hEF7: soft_out = 32'h02096F1B; // x = -4.1406, f(x) = 0.0159
    12'hEF8: soft_out = 32'h0211A538; // x = -4.1250, f(x) = 0.0162
    12'hEF9: soft_out = 32'h0219FC71; // x = -4.1094, f(x) = 0.0164
    12'hEFA: soft_out = 32'h02227549; // x = -4.0938, f(x) = 0.0167
    12'hEFB: soft_out = 32'h022B1048; // x = -4.0781, f(x) = 0.0169
    12'hEFC: soft_out = 32'h0233CDF9; // x = -4.0625, f(x) = 0.0172
    12'hEFD: soft_out = 32'h023CAEE7; // x = -4.0469, f(x) = 0.0175
    12'hEFE: soft_out = 32'h0245B3A0; // x = -4.0312, f(x) = 0.0178
    12'hEFF: soft_out = 32'h024EDCB5; // x = -4.0156, f(x) = 0.0180
    12'hF00: soft_out = 32'h02582AB7; // x = -4.0000, f(x) = 0.0183
    12'hF01: soft_out = 32'h02619E3C; // x = -3.9844, f(x) = 0.0186
    12'hF02: soft_out = 32'h026B37DC; // x = -3.9688, f(x) = 0.0189
    12'hF03: soft_out = 32'h0274F82F; // x = -3.9531, f(x) = 0.0192
    12'hF04: soft_out = 32'h027EDFD2; // x = -3.9375, f(x) = 0.0195
    12'hF05: soft_out = 32'h0288EF63; // x = -3.9219, f(x) = 0.0198
    12'hF06: soft_out = 32'h02932783; // x = -3.9062, f(x) = 0.0201
    12'hF07: soft_out = 32'h029D88D6; // x = -3.8906, f(x) = 0.0204
    12'hF08: soft_out = 32'h02A81401; // x = -3.8750, f(x) = 0.0208
    12'hF09: soft_out = 32'h02B2C9AE; // x = -3.8594, f(x) = 0.0211
    12'hF0A: soft_out = 32'h02BDAA88; // x = -3.8438, f(x) = 0.0214
    12'hF0B: soft_out = 32'h02C8B73D; // x = -3.8281, f(x) = 0.0218
    12'hF0C: soft_out = 32'h02D3F07E; // x = -3.8125, f(x) = 0.0221
    12'hF0D: soft_out = 32'h02DF56FD; // x = -3.7969, f(x) = 0.0224
    12'hF0E: soft_out = 32'h02EAEB73; // x = -3.7812, f(x) = 0.0228
    12'hF0F: soft_out = 32'h02F6AE97; // x = -3.7656, f(x) = 0.0232
    12'hF10: soft_out = 32'h0302A127; // x = -3.7500, f(x) = 0.0235
    12'hF11: soft_out = 32'h030EC3E1; // x = -3.7344, f(x) = 0.0239
    12'hF12: soft_out = 32'h031B1787; // x = -3.7188, f(x) = 0.0243
    12'hF13: soft_out = 32'h03279CDF; // x = -3.7031, f(x) = 0.0246
    12'hF14: soft_out = 32'h033454B1; // x = -3.6875, f(x) = 0.0250
    12'hF15: soft_out = 32'h03413FC9; // x = -3.6719, f(x) = 0.0254
    12'hF16: soft_out = 32'h034E5EF5; // x = -3.6562, f(x) = 0.0258
    12'hF17: soft_out = 32'h035BB307; // x = -3.6406, f(x) = 0.0262
    12'hF18: soft_out = 32'h03693CD5; // x = -3.6250, f(x) = 0.0266
    12'hF19: soft_out = 32'h0376FD37; // x = -3.6094, f(x) = 0.0271
    12'hF1A: soft_out = 32'h0384F508; // x = -3.5938, f(x) = 0.0275
    12'hF1B: soft_out = 32'h0393252A; // x = -3.5781, f(x) = 0.0279
    12'hF1C: soft_out = 32'h03A18E7E; // x = -3.5625, f(x) = 0.0284
    12'hF1D: soft_out = 32'h03B031EB; // x = -3.5469, f(x) = 0.0288
    12'hF1E: soft_out = 32'h03BF105C; // x = -3.5312, f(x) = 0.0293
    12'hF1F: soft_out = 32'h03CE2ABE; // x = -3.5156, f(x) = 0.0297
    12'hF20: soft_out = 32'h03DD8203; // x = -3.5000, f(x) = 0.0302
    12'hF21: soft_out = 32'h03ED1721; // x = -3.4844, f(x) = 0.0307
    12'hF22: soft_out = 32'h03FCEB10; // x = -3.4688, f(x) = 0.0312
    12'hF23: soft_out = 32'h040CFECE; // x = -3.4531, f(x) = 0.0316
    12'hF24: soft_out = 32'h041D535D; // x = -3.4375, f(x) = 0.0321
    12'hF25: soft_out = 32'h042DE9C1; // x = -3.4219, f(x) = 0.0327
    12'hF26: soft_out = 32'h043EC304; // x = -3.4062, f(x) = 0.0332
    12'hF27: soft_out = 32'h044FE034; // x = -3.3906, f(x) = 0.0337
    12'hF28: soft_out = 32'h04614262; // x = -3.3750, f(x) = 0.0342
    12'hF29: soft_out = 32'h0472EAA4; // x = -3.3594, f(x) = 0.0348
    12'hF2A: soft_out = 32'h0484DA16; // x = -3.3438, f(x) = 0.0353
    12'hF2B: soft_out = 32'h049711D5; // x = -3.3281, f(x) = 0.0359
    12'hF2C: soft_out = 32'h04A99306; // x = -3.3125, f(x) = 0.0364
    12'hF2D: soft_out = 32'h04BC5ED1; // x = -3.2969, f(x) = 0.0370
    12'hF2E: soft_out = 32'h04CF7662; // x = -3.2812, f(x) = 0.0376
    12'hF2F: soft_out = 32'h04E2DAEA; // x = -3.2656, f(x) = 0.0382
    12'hF30: soft_out = 32'h04F68DA1; // x = -3.2500, f(x) = 0.0388
    12'hF31: soft_out = 32'h050A8FC1; // x = -3.2344, f(x) = 0.0394
    12'hF32: soft_out = 32'h051EE28B; // x = -3.2188, f(x) = 0.0400
    12'hF33: soft_out = 32'h05338743; // x = -3.2031, f(x) = 0.0406
    12'hF34: soft_out = 32'h05487F34; // x = -3.1875, f(x) = 0.0413
    12'hF35: soft_out = 32'h055DCBAD; // x = -3.1719, f(x) = 0.0419
    12'hF36: soft_out = 32'h05736E04; // x = -3.1562, f(x) = 0.0426
    12'hF37: soft_out = 32'h05896792; // x = -3.1406, f(x) = 0.0433
    12'hF38: soft_out = 32'h059FB9B6; // x = -3.1250, f(x) = 0.0439
    12'hF39: soft_out = 32'h05B665D7; // x = -3.1094, f(x) = 0.0446
    12'hF3A: soft_out = 32'h05CD6D5F; // x = -3.0938, f(x) = 0.0453
    12'hF3B: soft_out = 32'h05E4D1BE; // x = -3.0781, f(x) = 0.0460
    12'hF3C: soft_out = 32'h05FC946B; // x = -3.0625, f(x) = 0.0468
    12'hF3D: soft_out = 32'h0614B6E1; // x = -3.0469, f(x) = 0.0475
    12'hF3E: soft_out = 32'h062D3AA4; // x = -3.0312, f(x) = 0.0483
    12'hF3F: soft_out = 32'h0646213A; // x = -3.0156, f(x) = 0.0490
    12'hF40: soft_out = 32'h065F6C33; // x = -3.0000, f(x) = 0.0498
    12'hF41: soft_out = 32'h06791D24; // x = -2.9844, f(x) = 0.0506
    12'hF42: soft_out = 32'h069335A6; // x = -2.9688, f(x) = 0.0514
    12'hF43: soft_out = 32'h06ADB75D; // x = -2.9531, f(x) = 0.0522
    12'hF44: soft_out = 32'h06C8A3F0; // x = -2.9375, f(x) = 0.0530
    12'hF45: soft_out = 32'h06E3FD0D; // x = -2.9219, f(x) = 0.0538
    12'hF46: soft_out = 32'h06FFC46B; // x = -2.9062, f(x) = 0.0547
    12'hF47: soft_out = 32'h071BFBC6; // x = -2.8906, f(x) = 0.0555
    12'hF48: soft_out = 32'h0738A4E1; // x = -2.8750, f(x) = 0.0564
    12'hF49: soft_out = 32'h0755C187; // x = -2.8594, f(x) = 0.0573
    12'hF4A: soft_out = 32'h0773538A; // x = -2.8438, f(x) = 0.0582
    12'hF4B: soft_out = 32'h07915CC2; // x = -2.8281, f(x) = 0.0591
    12'hF4C: soft_out = 32'h07AFDF11; // x = -2.8125, f(x) = 0.0601
    12'hF4D: soft_out = 32'h07CEDC5F; // x = -2.7969, f(x) = 0.0610
    12'hF4E: soft_out = 32'h07EE569B; // x = -2.7812, f(x) = 0.0620
    12'hF4F: soft_out = 32'h080E4FBD; // x = -2.7656, f(x) = 0.0629
    12'hF50: soft_out = 32'h082EC9C5; // x = -2.7500, f(x) = 0.0639
    12'hF51: soft_out = 32'h084FC6BA; // x = -2.7344, f(x) = 0.0649
    12'hF52: soft_out = 32'h087148AC; // x = -2.7188, f(x) = 0.0660
    12'hF53: soft_out = 32'h089351B3; // x = -2.7031, f(x) = 0.0670
    12'hF54: soft_out = 32'h08B5E3F0; // x = -2.6875, f(x) = 0.0681
    12'hF55: soft_out = 32'h08D9018C; // x = -2.6719, f(x) = 0.0691
    12'hF56: soft_out = 32'h08FCACB9; // x = -2.6562, f(x) = 0.0702
    12'hF57: soft_out = 32'h0920E7B2; // x = -2.6406, f(x) = 0.0713
    12'hF58: soft_out = 32'h0945B4BA; // x = -2.6250, f(x) = 0.0724
    12'hF59: soft_out = 32'h096B161E; // x = -2.6094, f(x) = 0.0736
    12'hF5A: soft_out = 32'h09910E34; // x = -2.5938, f(x) = 0.0747
    12'hF5B: soft_out = 32'h09B79F5B; // x = -2.5781, f(x) = 0.0759
    12'hF5C: soft_out = 32'h09DECBFE; // x = -2.5625, f(x) = 0.0771
    12'hF5D: soft_out = 32'h0A06968E; // x = -2.5469, f(x) = 0.0783
    12'hF5E: soft_out = 32'h0A2F0188; // x = -2.5312, f(x) = 0.0796
    12'hF5F: soft_out = 32'h0A580F73; // x = -2.5156, f(x) = 0.0808
    12'hF60: soft_out = 32'h0A81C2E0; // x = -2.5000, f(x) = 0.0821
    12'hF61: soft_out = 32'h0AAC1E6A; // x = -2.4844, f(x) = 0.0834
    12'hF62: soft_out = 32'h0AD724B7; // x = -2.4688, f(x) = 0.0847
    12'hF63: soft_out = 32'h0B02D877; // x = -2.4531, f(x) = 0.0860
    12'hF64: soft_out = 32'h0B2F3C66; // x = -2.4375, f(x) = 0.0874
    12'hF65: soft_out = 32'h0B5C5349; // x = -2.4219, f(x) = 0.0888
    12'hF66: soft_out = 32'h0B8A1FF3; // x = -2.4062, f(x) = 0.0902
    12'hF67: soft_out = 32'h0BB8A53F; // x = -2.3906, f(x) = 0.0916
    12'hF68: soft_out = 32'h0BE7E617; // x = -2.3750, f(x) = 0.0930
    12'hF69: soft_out = 32'h0C17E56E; // x = -2.3594, f(x) = 0.0945
    12'hF6A: soft_out = 32'h0C48A644; // x = -2.3438, f(x) = 0.0960
    12'hF6B: soft_out = 32'h0C7A2BA6; // x = -2.3281, f(x) = 0.0975
    12'hF6C: soft_out = 32'h0CAC78AB; // x = -2.3125, f(x) = 0.0990
    12'hF6D: soft_out = 32'h0CDF907A; // x = -2.2969, f(x) = 0.1006
    12'hF6E: soft_out = 32'h0D137642; // x = -2.2812, f(x) = 0.1022
    12'hF6F: soft_out = 32'h0D482D43; // x = -2.2656, f(x) = 0.1038
    12'hF70: soft_out = 32'h0D7DB8C7; // x = -2.2500, f(x) = 0.1054
    12'hF71: soft_out = 32'h0DB41C29; // x = -2.2344, f(x) = 0.1071
    12'hF72: soft_out = 32'h0DEB5ACD; // x = -2.2188, f(x) = 0.1087
    12'hF73: soft_out = 32'h0E237828; // x = -2.2031, f(x) = 0.1105
    12'hF74: soft_out = 32'h0E5C77BC; // x = -2.1875, f(x) = 0.1122
    12'hF75: soft_out = 32'h0E965D18; // x = -2.1719, f(x) = 0.1140
    12'hF76: soft_out = 32'h0ED12BDC; // x = -2.1562, f(x) = 0.1158
    12'hF77: soft_out = 32'h0F0CE7B3; // x = -2.1406, f(x) = 0.1176
    12'hF78: soft_out = 32'h0F49945A; // x = -2.1250, f(x) = 0.1194
    12'hF79: soft_out = 32'h0F87359C; // x = -2.1094, f(x) = 0.1213
    12'hF7A: soft_out = 32'h0FC5CF53; // x = -2.0938, f(x) = 0.1232
    12'hF7B: soft_out = 32'h10056567; // x = -2.0781, f(x) = 0.1252
    12'hF7C: soft_out = 32'h1045FBD4; // x = -2.0625, f(x) = 0.1271
    12'hF7D: soft_out = 32'h108796A1; // x = -2.0469, f(x) = 0.1291
    12'hF7E: soft_out = 32'h10CA39E9; // x = -2.0312, f(x) = 0.1312
    12'hF7F: soft_out = 32'h110DE9D6; // x = -2.0156, f(x) = 0.1332
    12'hF80: soft_out = 32'h1152AAA4; // x = -2.0000, f(x) = 0.1353
    12'hF81: soft_out = 32'h1198809D; // x = -1.9844, f(x) = 0.1375
    12'hF82: soft_out = 32'h11DF7020; // x = -1.9688, f(x) = 0.1396
    12'hF83: soft_out = 32'h12277D9B; // x = -1.9531, f(x) = 0.1418
    12'hF84: soft_out = 32'h1270AD90; // x = -1.9375, f(x) = 0.1441
    12'hF85: soft_out = 32'h12BB0491; // x = -1.9219, f(x) = 0.1463
    12'hF86: soft_out = 32'h13068744; // x = -1.9062, f(x) = 0.1486
    12'hF87: soft_out = 32'h13533A61; // x = -1.8906, f(x) = 0.1510
    12'hF88: soft_out = 32'h13A122B4; // x = -1.8750, f(x) = 0.1534
    12'hF89: soft_out = 32'h13F0451A; // x = -1.8594, f(x) = 0.1558
    12'hF8A: soft_out = 32'h1440A686; // x = -1.8438, f(x) = 0.1582
    12'hF8B: soft_out = 32'h14924BFE; // x = -1.8281, f(x) = 0.1607
    12'hF8C: soft_out = 32'h14E53A9D; // x = -1.8125, f(x) = 0.1632
    12'hF8D: soft_out = 32'h15397791; // x = -1.7969, f(x) = 0.1658
    12'hF8E: soft_out = 32'h158F081E; // x = -1.7812, f(x) = 0.1684
    12'hF8F: soft_out = 32'h15E5F19E; // x = -1.7656, f(x) = 0.1711
    12'hF90: soft_out = 32'h163E397E; // x = -1.7500, f(x) = 0.1738
    12'hF91: soft_out = 32'h1697E544; // x = -1.7344, f(x) = 0.1765
    12'hF92: soft_out = 32'h16F2FA8A; // x = -1.7188, f(x) = 0.1793
    12'hF93: soft_out = 32'h174F7F02; // x = -1.7031, f(x) = 0.1821
    12'hF94: soft_out = 32'h17AD7873; // x = -1.6875, f(x) = 0.1850
    12'hF95: soft_out = 32'h180CECBF; // x = -1.6719, f(x) = 0.1879
    12'hF96: soft_out = 32'h186DE1DB; // x = -1.6562, f(x) = 0.1909
    12'hF97: soft_out = 32'h18D05DD7; // x = -1.6406, f(x) = 0.1939
    12'hF98: soft_out = 32'h193466DB; // x = -1.6250, f(x) = 0.1969
    12'hF99: soft_out = 32'h199A0327; // x = -1.6094, f(x) = 0.2000
    12'hF9A: soft_out = 32'h1A013916; // x = -1.5938, f(x) = 0.2032
    12'hF9B: soft_out = 32'h1A6A0F1B; // x = -1.5781, f(x) = 0.2064
    12'hF9C: soft_out = 32'h1AD48BC2; // x = -1.5625, f(x) = 0.2096
    12'hF9D: soft_out = 32'h1B40B5B5; // x = -1.5469, f(x) = 0.2129
    12'hF9E: soft_out = 32'h1BAE93B5; // x = -1.5312, f(x) = 0.2163
    12'hF9F: soft_out = 32'h1C1E2CA1; // x = -1.5156, f(x) = 0.2197
    12'hFA0: soft_out = 32'h1C8F8772; // x = -1.5000, f(x) = 0.2231
    12'hFA1: soft_out = 32'h1D02AB3E; // x = -1.4844, f(x) = 0.2266
    12'hFA2: soft_out = 32'h1D779F37; // x = -1.4688, f(x) = 0.2302
    12'hFA3: soft_out = 32'h1DEE6AAD; // x = -1.4531, f(x) = 0.2338
    12'hFA4: soft_out = 32'h1E67150B; // x = -1.4375, f(x) = 0.2375
    12'hFA5: soft_out = 32'h1EE1A5DD; // x = -1.4219, f(x) = 0.2413
    12'hFA6: soft_out = 32'h1F5E24CD; // x = -1.4062, f(x) = 0.2451
    12'hFA7: soft_out = 32'h1FDC99A1; // x = -1.3906, f(x) = 0.2489
    12'hFA8: soft_out = 32'h205D0C42; // x = -1.3750, f(x) = 0.2528
    12'hFA9: soft_out = 32'h20DF84B6; // x = -1.3594, f(x) = 0.2568
    12'hFAA: soft_out = 32'h21640B25; // x = -1.3438, f(x) = 0.2609
    12'hFAB: soft_out = 32'h21EAA7D7; // x = -1.3281, f(x) = 0.2650
    12'hFAC: soft_out = 32'h22736337; // x = -1.3125, f(x) = 0.2691
    12'hFAD: soft_out = 32'h22FE45D0; // x = -1.2969, f(x) = 0.2734
    12'hFAE: soft_out = 32'h238B5850; // x = -1.2812, f(x) = 0.2777
    12'hFAF: soft_out = 32'h241AA388; // x = -1.2656, f(x) = 0.2821
    12'hFB0: soft_out = 32'h24AC306E; // x = -1.2500, f(x) = 0.2865
    12'hFB1: soft_out = 32'h2540081A; // x = -1.2344, f(x) = 0.2910
    12'hFB2: soft_out = 32'h25D633CA; // x = -1.2188, f(x) = 0.2956
    12'hFB3: soft_out = 32'h266EBCE0; // x = -1.2031, f(x) = 0.3003
    12'hFB4: soft_out = 32'h2709ACE5; // x = -1.1875, f(x) = 0.3050
    12'hFB5: soft_out = 32'h27A70D88; // x = -1.1719, f(x) = 0.3098
    12'hFB6: soft_out = 32'h2846E89F; // x = -1.1562, f(x) = 0.3147
    12'hFB7: soft_out = 32'h28E94828; // x = -1.1406, f(x) = 0.3196
    12'hFB8: soft_out = 32'h298E3649; // x = -1.1250, f(x) = 0.3247
    12'hFB9: soft_out = 32'h2A35BD51; // x = -1.1094, f(x) = 0.3298
    12'hFBA: soft_out = 32'h2ADFE7B8; // x = -1.0938, f(x) = 0.3350
    12'hFBB: soft_out = 32'h2B8CC021; // x = -1.0781, f(x) = 0.3402
    12'hFBC: soft_out = 32'h2C3C515A; // x = -1.0625, f(x) = 0.3456
    12'hFBD: soft_out = 32'h2CEEA65C; // x = -1.0469, f(x) = 0.3510
    12'hFBE: soft_out = 32'h2DA3CA4B; // x = -1.0312, f(x) = 0.3566
    12'hFBF: soft_out = 32'h2E5BC87C; // x = -1.0156, f(x) = 0.3622
    12'hFC0: soft_out = 32'h2F16AC6C; // x = -1.0000, f(x) = 0.3679
    12'hFC1: soft_out = 32'h2FD481CC; // x = -0.9844, f(x) = 0.3737
    12'hFC2: soft_out = 32'h30955477; // x = -0.9688, f(x) = 0.3796
    12'hFC3: soft_out = 32'h3159307C; // x = -0.9531, f(x) = 0.3855
    12'hFC4: soft_out = 32'h32202218; // x = -0.9375, f(x) = 0.3916
    12'hFC5: soft_out = 32'h32EA35BA; // x = -0.9219, f(x) = 0.3978
    12'hFC6: soft_out = 32'h33B77804; // x = -0.9062, f(x) = 0.4040
    12'hFC7: soft_out = 32'h3487F5C9; // x = -0.8906, f(x) = 0.4104
    12'hFC8: soft_out = 32'h355BBC13; // x = -0.8750, f(x) = 0.4169
    12'hFC9: soft_out = 32'h3632D81C; // x = -0.8594, f(x) = 0.4234
    12'hFCA: soft_out = 32'h370D5758; // x = -0.8438, f(x) = 0.4301
    12'hFCB: soft_out = 32'h37EB476D; // x = -0.8281, f(x) = 0.4369
    12'hFCC: soft_out = 32'h38CCB63C; // x = -0.8125, f(x) = 0.4437
    12'hFCD: soft_out = 32'h39B1B1DB; // x = -0.7969, f(x) = 0.4507
    12'hFCE: soft_out = 32'h3A9A489A; // x = -0.7812, f(x) = 0.4578
    12'hFCF: soft_out = 32'h3B868902; // x = -0.7656, f(x) = 0.4650
    12'hFD0: soft_out = 32'h3C7681D8; // x = -0.7500, f(x) = 0.4724
    12'hFD1: soft_out = 32'h3D6A421B; // x = -0.7344, f(x) = 0.4798
    12'hFD2: soft_out = 32'h3E61D907; // x = -0.7188, f(x) = 0.4874
    12'hFD3: soft_out = 32'h3F5D5616; // x = -0.7031, f(x) = 0.4950
    12'hFD4: soft_out = 32'h405CC8FF; // x = -0.6875, f(x) = 0.5028
    12'hFD5: soft_out = 32'h416041BB; // x = -0.6719, f(x) = 0.5108
    12'hFD6: soft_out = 32'h4267D080; // x = -0.6562, f(x) = 0.5188
    12'hFD7: soft_out = 32'h437385C8; // x = -0.6406, f(x) = 0.5270
    12'hFD8: soft_out = 32'h4483724D; // x = -0.6250, f(x) = 0.5353
    12'hFD9: soft_out = 32'h4597A710; // x = -0.6094, f(x) = 0.5437
    12'hFDA: soft_out = 32'h46B03552; // x = -0.5938, f(x) = 0.5523
    12'hFDB: soft_out = 32'h47CD2E9E; // x = -0.5781, f(x) = 0.5609
    12'hFDC: soft_out = 32'h48EEA4C3; // x = -0.5625, f(x) = 0.5698
    12'hFDD: soft_out = 32'h4A14A9D8; // x = -0.5469, f(x) = 0.5788
    12'hFDE: soft_out = 32'h4B3F503E; // x = -0.5312, f(x) = 0.5879
    12'hFDF: soft_out = 32'h4C6EAA9F; // x = -0.5156, f(x) = 0.5971
    12'hFE0: soft_out = 32'h4DA2CBF2; // x = -0.5000, f(x) = 0.6065
    12'hFE1: soft_out = 32'h4EDBC777; // x = -0.4844, f(x) = 0.6161
    12'hFE2: soft_out = 32'h5019B0C0; // x = -0.4688, f(x) = 0.6258
    12'hFE3: soft_out = 32'h515C9BAA; // x = -0.4531, f(x) = 0.6356
    12'hFE4: soft_out = 32'h52A49C65; // x = -0.4375, f(x) = 0.6456
    12'hFE5: soft_out = 32'h53F1C770; // x = -0.4219, f(x) = 0.6558
    12'hFE6: soft_out = 32'h5544319F; // x = -0.4062, f(x) = 0.6661
    12'hFE7: soft_out = 32'h569BF018; // x = -0.3906, f(x) = 0.6766
    12'hFE8: soft_out = 32'h57F91858; // x = -0.3750, f(x) = 0.6873
    12'hFE9: soft_out = 32'h595BC030; // x = -0.3594, f(x) = 0.6981
    12'hFEA: soft_out = 32'h5AC3FDCB; // x = -0.3438, f(x) = 0.7091
    12'hFEB: soft_out = 32'h5C31E7AF; // x = -0.3281, f(x) = 0.7203
    12'hFEC: soft_out = 32'h5DA594B8; // x = -0.3125, f(x) = 0.7316
    12'hFED: soft_out = 32'h5F1F1C22; // x = -0.2969, f(x) = 0.7431
    12'hFEE: soft_out = 32'h609E9586; // x = -0.2812, f(x) = 0.7548
    12'hFEF: soft_out = 32'h622418DC; // x = -0.2656, f(x) = 0.7667
    12'hFF0: soft_out = 32'h63AFBE7B; // x = -0.2500, f(x) = 0.7788
    12'hFF1: soft_out = 32'h65419F1E; // x = -0.2344, f(x) = 0.7911
    12'hFF2: soft_out = 32'h66D9D3E4; // x = -0.2188, f(x) = 0.8035
    12'hFF3: soft_out = 32'h6878764F; // x = -0.2031, f(x) = 0.8162
    12'hFF4: soft_out = 32'h6A1DA04B; // x = -0.1875, f(x) = 0.8290
    12'hFF5: soft_out = 32'h6BC96C2A; // x = -0.1719, f(x) = 0.8421
    12'hFF6: soft_out = 32'h6D7BF4A8; // x = -0.1562, f(x) = 0.8553
    12'hFF7: soft_out = 32'h6F3554EE; // x = -0.1406, f(x) = 0.8688
    12'hFF8: soft_out = 32'h70F5A894; // x = -0.1250, f(x) = 0.8825
    12'hFF9: soft_out = 32'h72BD0B9D; // x = -0.1094, f(x) = 0.8964
    12'hFFA: soft_out = 32'h748B9A80; // x = -0.0938, f(x) = 0.9105
    12'hFFB: soft_out = 32'h76617227; // x = -0.0781, f(x) = 0.9248
    12'hFFC: soft_out = 32'h783EAFEF; // x = -0.0625, f(x) = 0.9394
    12'hFFD: soft_out = 32'h7A2371AC; // x = -0.0469, f(x) = 0.9542
    12'hFFE: soft_out = 32'h7C0FD5AA; // x = -0.0312, f(x) = 0.9692
    12'hFFF: soft_out = 32'h7E03FAB0; // x = -0.0156, f(x) = 0.9845
    default: soft_out = 32'h0; 
  endcase
end

//------------------------------------------------------------------------
// FSM
//------------------------------------------------------------------------

localparam IDLE    = 2'd0;
localparam EXP     = 2'd1;
localparam RECIP   = 2'd2;
localparam SOFTMAX = 2'd3;

localparam Exponential = 2'd0;
localparam Reciprocal  = 2'd1;
localparam Softmax     = 2'd2;

reg [2:0] curr_state, next_state;

always@ ( posedge clk ) begin
    if ( reset ) begin
      curr_state <= IDLE;
    end
    else begin
      curr_state <= next_state;
    end
end

always@ (*) begin
    next_state = curr_state;
    case ( curr_state )
      IDLE  : begin
        if ( cmd_valid ) begin
          case ( cmd_payload_function_id[9:3] )
            Exponential: next_state = EXP;
            Reciprocal : next_state = RECIP;
            Softmax    : next_state = SOFTMAX;
            default    : next_state = IDLE;
          endcase
        end
      end
      EXP    : next_state = ( rsp_ready ) ? IDLE : EXP;
      RECIP  : next_state = ( rsp_ready ) ? IDLE : RECIP;
      SOFTMAX: next_state = ( rsp_ready ) ? IDLE : SOFTMAX;
      default: next_state = IDLE;
    endcase
end


always@ (*) begin
    cmd_ready             = 1'b0;
    rsp_valid             = 1'b0;
    rsp_payload_outputs_0 = 32'd0;
    case ( curr_state )
      IDLE: begin
        cmd_ready = 1'b1;
        rsp_valid = 1'b0;
        rsp_payload_outputs_0 = 32'd0;
      end
      EXP: begin
        cmd_ready = 1'b0;
        rsp_valid = 1'b1;
        rsp_payload_outputs_0 = exp_out;
      end
      RECIP: begin
        cmd_ready = 1'b0;
        rsp_valid = 1'b1;
        rsp_payload_outputs_0 = recip_out;
      end      
      SOFTMAX: begin
        cmd_ready = 1'b0;
        rsp_valid = 1'b1;
        rsp_payload_outputs_0 = soft_out;
      end
    endcase
end

endmodule
